`timescale 1ns / 1ps
`include "modulator_signals.vh"

module baseband_dsp_tb;

    reg data_in;
    reg data_clk;
    reg dsp_clk;
    reg rst_n_data;
    reg rst_n_dsp;
    reg msg_in;
    reg rw;
    reg [9:0] mem_addr;
    reg [7:0] coeff_in; 
    reg enable;
    reg [3:0] sample_rate;
    reg mapping;
    wire mem_read_out;
    wire [9:0] I_out;
    wire [9:0] Q_out;

    baseband_dsp DUT(
        .data_in(data_in),
        .data_clk(data_clk),
        .dsp_clk(dsp_clk),
        .rst_n_data(rst_n_data),
        .rst_n_dsp(rst_n_dsp),
        .msg_in(msg_in),
        .rw(rw),
        .mem_addr(mem_addr),
        .coeff_in(coeff_in),
        .mem_read_out(mem_read_out),
        .I_out(I_out),
	    .Q_out(Q_out)
    );
	
	// Datastream variables
	reg [7:0] Icoeff [0:70];
	reg [7:0] Qcoeff [0:70];
	reg [779:0] datastream;
	reg [9:0] I_filtered_10b[0:1733];
	reg [9:0] Q_filtered_10b[0:1733];
	reg [11:0] I_filtered_12b[0:63]; //11
	reg [11:0] Q_filtered_12b[0:63]; //11
	
    always #8.333 data_clk = ~data_clk;
    always #3.846 dsp_clk = ~dsp_clk;
    
    reg [8*39:0] testcase;
    integer i;
	
    initial begin
        testcase = "Initializing";
        data_clk <= 1'b0;
        dsp_clk <= 1'b0;
        rst_n_data <= 1'b0;
        rst_n_dsp <= 1'b0;
		sample_rate <= 4'd13;
        data_in <= 1'b0; 
        enable <= 1'b0;

		repeat(2) @(posedge data_clk);
		rst_n_data <= 1'b1;
        enable <= 1'b1;
		@(posedge data_clk);

        @(posedge dsp_clk)
        rst_n_dsp <= 1'b1;
        @(posedge dsp_clk)

        // Write I coefficients to memory
        @(negedge dsp_clk);
		for (i=0; i<=70; i=i+1) begin
			msg_in <= 1'b1;
			rw <= 1'b1;
			mem_addr  <= i + 128;
			coeff_in  <= Icoeff[i];
			@(negedge dsp_clk);	 
		end

		// Write Q coefficients to memory
		for (i=0; i<=70; i = i+1) begin
			msg_in <= 1'b1;
			rw <= 1'b1;
			mem_addr  <= i + 256;
			coeff_in  <= Qcoeff[i];
			@(negedge dsp_clk);	 
		end
		msg_in <= 1'b0;

        testcase = "Coeff_Read";
        repeat(3) @(posedge dsp_clk);
        // Test reading coeff I memory
		// coeff_read_out should set to 0xFD
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr  <= 133; // This is addr of 5th I coeff: oxFD
		repeat(2) @(posedge dsp_clk);
		msg_in <= 1'b0;

		repeat(3) @(posedge dsp_clk);
		// Test reading coeff Q memory
		// coeff_read_out should set to 0x02
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr  <= 266; 
		repeat(3) @(posedge dsp_clk);
		msg_in <= 1'b0;

		// flush the pipeline
		repeat(5) @(posedge dsp_clk);

        // Send in datastream with 12 bit header
        testcase <= "Datastream";    
        @(negedge data_clk);
        for (i=779; i>=0; i=i-1) begin
            data_in <= datastream[i]; 
            @(negedge data_clk);
        end

        repeat(3) @(posedge dsp_clk);
        // Test reading I output memory
		// Should read 10th output: 0x00 or 0x05F idk
        testcase <= "Output_read"; 
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr <= 512;
		// Read last 4 LSBs
		repeat(1) @(posedge dsp_clk);
		mem_addr  <= 513;
		repeat(3) @(posedge dsp_clk);

		// Test reading I output memory
		// Should read 10th output: 0x090 or 0x082 or 0xFF6 idk
        testcase <= "Output_read"; 
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr <= 532;
		// Read last 4 LSBs
		repeat(1) @(posedge dsp_clk);
		mem_addr  <= 533;
		repeat(3) @(posedge dsp_clk);

        // Write compare outputs function and log file
        $finish;
    end

initial begin
    // I filter coefficients
    Icoeff[0] = 00;
    Icoeff[1] = 00;
    Icoeff[2] = FF;
    Icoeff[3] = FE;
    Icoeff[4] = FE;
    Icoeff[5] = FD;
    Icoeff[6] = FE;
    Icoeff[7] = FE;
    Icoeff[8] = FF;
    Icoeff[9] = 00;
    Icoeff[10] = 02;
    Icoeff[11] = 03;
    Icoeff[12] = 03;
    Icoeff[13] = 03;
    Icoeff[14] = 02;
    Icoeff[15] = 01;
    Icoeff[16] = FE;
    Icoeff[17] = FB;
    Icoeff[18] = F8;
    Icoeff[19] = F5;
    Icoeff[20] = F3;
    Icoeff[21] = F3;
    Icoeff[22] = F4;
    Icoeff[23] = F7;
    Icoeff[24] = FE;
    Icoeff[25] = 07;
    Icoeff[26] = 12;
    Icoeff[27] = 20;
    Icoeff[28] = 30;
    Icoeff[29] = 40;
    Icoeff[30] = 51;
    Icoeff[31] = 60;
    Icoeff[32] = 6D;
    Icoeff[33] = 77;
    Icoeff[34] = 7D;
    Icoeff[35] = 7F;
    Icoeff[36] = 7D;
    Icoeff[37] = 77;
    Icoeff[38] = 6D;
    Icoeff[39] = 60;
    Icoeff[40] = 51;
    Icoeff[41] = 40;
    Icoeff[42] = 30;
    Icoeff[43] = 20;
    Icoeff[44] = 12;
    Icoeff[45] = 07;
    Icoeff[46] = FE;
    Icoeff[47] = F7;
    Icoeff[48] = F4;
    Icoeff[49] = F3;
    Icoeff[50] = F3;
    Icoeff[51] = F5;
    Icoeff[52] = F8;
    Icoeff[53] = FB;
    Icoeff[54] = FE;
    Icoeff[55] = 01;
    Icoeff[56] = 02;
    Icoeff[57] = 03;
    Icoeff[58] = 03;
    Icoeff[59] = 03;
    Icoeff[60] = 02;
    Icoeff[61] = 00;
    Icoeff[62] = FF;
    Icoeff[63] = FE;
    Icoeff[64] = FE;
    Icoeff[65] = FD;
    Icoeff[66] = FE;
    Icoeff[67] = FE;
    Icoeff[68] = FF;
    Icoeff[69] = 00;
    Icoeff[70] = 00;


// Q filter coefficients
    Qcoeff[0] = 00;
    Qcoeff[1] = 00;
    Qcoeff[2] = FF;
    Qcoeff[3] = FE;
    Qcoeff[4] = FE;
    Qcoeff[5] = FD;
    Qcoeff[6] = FE;
    Qcoeff[7] = FE;
    Qcoeff[8] = FF;
    Qcoeff[9] = 00;
    Qcoeff[10] = 02;
    Qcoeff[11] = 03;
    Qcoeff[12] = 03;
    Qcoeff[13] = 03;
    Qcoeff[14] = 02;
    Qcoeff[15] = 01;
    Qcoeff[16] = FE;
    Qcoeff[17] = FB;
    Qcoeff[18] = F9;
    Qcoeff[19] = F6;
    Qcoeff[20] = F4;
    Qcoeff[21] = F4;
    Qcoeff[22] = F5;
    Qcoeff[23] = F8;
    Qcoeff[24] = FE;
    Qcoeff[25] = 06;
    Qcoeff[26] = 10;
    Qcoeff[27] = 1D;
    Qcoeff[28] = 2B;
    Qcoeff[29] = 3A;
    Qcoeff[30] = 49;
    Qcoeff[31] = 56;
    Qcoeff[32] = 62;
    Qcoeff[33] = 6B;
    Qcoeff[34] = 71;
    Qcoeff[35] = 72;
    Qcoeff[36] = 71;
    Qcoeff[37] = 6B;
    Qcoeff[38] = 62;
    Qcoeff[39] = 56;
    Qcoeff[40] = 49;
    Qcoeff[41] = 3A;
    Qcoeff[42] = 2B;
    Qcoeff[43] = 1D;
    Qcoeff[44] = 10;
    Qcoeff[45] = 06;
    Qcoeff[46] = FE;
    Qcoeff[47] = F8;
    Qcoeff[48] = F5;
    Qcoeff[49] = F4;
    Qcoeff[50] = F4;
    Qcoeff[51] = F6;
    Qcoeff[52] = F9;
    Qcoeff[53] = FB;
    Qcoeff[54] = FE;
    Qcoeff[55] = 01;
    Qcoeff[56] = 02;
    Qcoeff[57] = 03;
    Qcoeff[58] = 03;
    Qcoeff[59] = 03;
    Qcoeff[60] = 02;
    Qcoeff[61] = 00;
    Qcoeff[62] = FF;
    Qcoeff[63] = FE;
    Qcoeff[64] = FE;
    Qcoeff[65] = FD;
    Qcoeff[66] = FE;
    Qcoeff[67] = FE;
    Qcoeff[68] = FF;
    Qcoeff[69] = 00;
    Qcoeff[70] = 00;


// Transmit Datastream with header
    [779:768] datastream = B38;
    [767:752] datastream = D196;
    [751:736] datastream = 7592;
    [735:720] datastream = FAE7;
    [719:704] datastream = 8104;
    [703:688] datastream = 35D3;
    [687:672] datastream = 6897;
    [671:656] datastream = 9BF2;
    [655:640] datastream = A590;
    [639:624] datastream = 451B;
    [623:608] datastream = E113;
    [607:592] datastream = 15AC;
    [591:576] datastream = CB73;
    [575:560] datastream = DEBF;
    [559:544] datastream = 0193;
    [543:528] datastream = 6465;
    [527:512] datastream = 02F3;
    [511:496] datastream = 9786;
    [495:480] datastream = 4A79;
    [479:464] datastream = 6B6F;
    [463:448] datastream = 2E55;
    [447:432] datastream = CDA6;
    [431:416] datastream = 8028;
    [415:400] datastream = 5FE6;
    [399:384] datastream = 80E7;
    [383:368] datastream = FE45;
    [367:352] datastream = 8CF6;
    [351:336] datastream = C49A;
    [335:320] datastream = 4E25;
    [319:304] datastream = F8C8;
    [303:288] datastream = 0985;
    [287:272] datastream = FC5F;
    [271:256] datastream = 23B5;
    [255:240] datastream = 94F7;
    [239:224] datastream = B931;
    [223:208] datastream = E1FA;
    [207:192] datastream = 6604;
    [191:176] datastream = CB9A;
    [175:160] datastream = EA5C;
    [159:144] datastream = 2DE4;
    [143:128] datastream = F7BA;
    [127:112] datastream = 962F;
    [111:96] datastream = 329D;
    [95:80] datastream = 7727;
    [79:64] datastream = 9533;
    [63:48] datastream = 2149;
    [47:32] datastream = 386A;
    [31:16] datastream = E179;
    [15:0] datastream = AA26;


// I Channel 10b Expected output
    I_filtered_10b[1733] = 000;
    I_filtered_10b[1732] = 000;
    I_filtered_10b[1731] = 000;
    I_filtered_10b[1730] = 000;
    I_filtered_10b[1729] = 000;
    I_filtered_10b[1728] = 000;
    I_filtered_10b[1727] = 000;
    I_filtered_10b[1726] = 000;
    I_filtered_10b[1725] = 000;
    I_filtered_10b[1724] = 000;
    I_filtered_10b[1723] = 000;
    I_filtered_10b[1722] = 000;
    I_filtered_10b[1721] = 000;
    I_filtered_10b[1720] = 000;
    I_filtered_10b[1719] = 000;
    I_filtered_10b[1718] = 000;
    I_filtered_10b[1717] = 000;
    I_filtered_10b[1716] = 001;
    I_filtered_10b[1715] = 000;
    I_filtered_10b[1714] = 000;
    I_filtered_10b[1713] = 000;
    I_filtered_10b[1712] = 000;
    I_filtered_10b[1711] = 000;
    I_filtered_10b[1710] = 3FF;
    I_filtered_10b[1709] = 3FF;
    I_filtered_10b[1708] = 3FF;
    I_filtered_10b[1707] = 000;
    I_filtered_10b[1706] = 001;
    I_filtered_10b[1705] = 004;
    I_filtered_10b[1704] = 005;
    I_filtered_10b[1703] = 007;
    I_filtered_10b[1702] = 006;
    I_filtered_10b[1701] = 007;
    I_filtered_10b[1700] = 005;
    I_filtered_10b[1699] = 003;
    I_filtered_10b[1698] = 3FF;
    I_filtered_10b[1697] = 3FB;
    I_filtered_10b[1696] = 3F9;
    I_filtered_10b[1695] = 3F6;
    I_filtered_10b[1694] = 3F5;
    I_filtered_10b[1693] = 3F3;
    I_filtered_10b[1692] = 3F5;
    I_filtered_10b[1691] = 3F6;
    I_filtered_10b[1690] = 3F8;
    I_filtered_10b[1689] = 3FA;
    I_filtered_10b[1688] = 3FB;
    I_filtered_10b[1687] = 3F8;
    I_filtered_10b[1686] = 3F5;
    I_filtered_10b[1685] = 3EF;
    I_filtered_10b[1684] = 3E4;
    I_filtered_10b[1683] = 3D6;
    I_filtered_10b[1682] = 3C6;
    I_filtered_10b[1681] = 3B2;
    I_filtered_10b[1680] = 39C;
    I_filtered_10b[1679] = 386;
    I_filtered_10b[1678] = 36F;
    I_filtered_10b[1677] = 35A;
    I_filtered_10b[1676] = 348;
    I_filtered_10b[1675] = 33B;
    I_filtered_10b[1674] = 332;
    I_filtered_10b[1673] = 32E;
    I_filtered_10b[1672] = 32F;
    I_filtered_10b[1671] = 334;
    I_filtered_10b[1670] = 33E;
    I_filtered_10b[1669] = 34C;
    I_filtered_10b[1668] = 35B;
    I_filtered_10b[1667] = 36C;
    I_filtered_10b[1666] = 37C;
    I_filtered_10b[1665] = 38C;
    I_filtered_10b[1664] = 399;
    I_filtered_10b[1663] = 3A4;
    I_filtered_10b[1662] = 3AC;
    I_filtered_10b[1661] = 3B5;
    I_filtered_10b[1660] = 3B9;
    I_filtered_10b[1659] = 3BC;
    I_filtered_10b[1658] = 3BF;
    I_filtered_10b[1657] = 3C1;
    I_filtered_10b[1656] = 3C3;
    I_filtered_10b[1655] = 3C5;
    I_filtered_10b[1654] = 3C7;
    I_filtered_10b[1653] = 3C8;
    I_filtered_10b[1652] = 3CD;
    I_filtered_10b[1651] = 3D0;
    I_filtered_10b[1650] = 3D5;
    I_filtered_10b[1649] = 3D9;
    I_filtered_10b[1648] = 3E0;
    I_filtered_10b[1647] = 3E6;
    I_filtered_10b[1646] = 3ED;
    I_filtered_10b[1645] = 3F3;
    I_filtered_10b[1644] = 3F6;
    I_filtered_10b[1643] = 3FC;
    I_filtered_10b[1642] = 3FE;
    I_filtered_10b[1641] = 002;
    I_filtered_10b[1640] = 003;
    I_filtered_10b[1639] = 005;
    I_filtered_10b[1638] = 008;
    I_filtered_10b[1637] = 00A;
    I_filtered_10b[1636] = 00C;
    I_filtered_10b[1635] = 010;
    I_filtered_10b[1634] = 014;
    I_filtered_10b[1633] = 017;
    I_filtered_10b[1632] = 01F;
    I_filtered_10b[1631] = 027;
    I_filtered_10b[1630] = 032;
    I_filtered_10b[1629] = 03E;
    I_filtered_10b[1628] = 04E;
    I_filtered_10b[1627] = 05D;
    I_filtered_10b[1626] = 06E;
    I_filtered_10b[1625] = 07E;
    I_filtered_10b[1624] = 08C;
    I_filtered_10b[1623] = 097;
    I_filtered_10b[1622] = 09D;
    I_filtered_10b[1621] = 09F;
    I_filtered_10b[1620] = 09B;
    I_filtered_10b[1619] = 092;
    I_filtered_10b[1618] = 083;
    I_filtered_10b[1617] = 071;
    I_filtered_10b[1616] = 05C;
    I_filtered_10b[1615] = 043;
    I_filtered_10b[1614] = 02C;
    I_filtered_10b[1613] = 015;
    I_filtered_10b[1612] = 000;
    I_filtered_10b[1611] = 3F1;
    I_filtered_10b[1610] = 3E3;
    I_filtered_10b[1609] = 3D9;
    I_filtered_10b[1608] = 3D4;
    I_filtered_10b[1607] = 3D3;
    I_filtered_10b[1606] = 3D3;
    I_filtered_10b[1605] = 3D6;
    I_filtered_10b[1604] = 3DA;
    I_filtered_10b[1603] = 3DE;
    I_filtered_10b[1602] = 3E1;
    I_filtered_10b[1601] = 3E3;
    I_filtered_10b[1600] = 3E4;
    I_filtered_10b[1599] = 3E3;
    I_filtered_10b[1598] = 3E3;
    I_filtered_10b[1597] = 3E2;
    I_filtered_10b[1596] = 3E2;
    I_filtered_10b[1595] = 3E0;
    I_filtered_10b[1594] = 3E2;
    I_filtered_10b[1593] = 3E5;
    I_filtered_10b[1592] = 3E9;
    I_filtered_10b[1591] = 3ED;
    I_filtered_10b[1590] = 3F4;
    I_filtered_10b[1589] = 3FC;
    I_filtered_10b[1588] = 002;
    I_filtered_10b[1587] = 009;
    I_filtered_10b[1586] = 00F;
    I_filtered_10b[1585] = 012;
    I_filtered_10b[1584] = 015;
    I_filtered_10b[1583] = 018;
    I_filtered_10b[1582] = 01A;
    I_filtered_10b[1581] = 01A;
    I_filtered_10b[1580] = 01E;
    I_filtered_10b[1579] = 021;
    I_filtered_10b[1578] = 026;
    I_filtered_10b[1577] = 02C;
    I_filtered_10b[1576] = 035;
    I_filtered_10b[1575] = 040;
    I_filtered_10b[1574] = 04A;
    I_filtered_10b[1573] = 055;
    I_filtered_10b[1572] = 05D;
    I_filtered_10b[1571] = 064;
    I_filtered_10b[1570] = 066;
    I_filtered_10b[1569] = 065;
    I_filtered_10b[1568] = 05F;
    I_filtered_10b[1567] = 054;
    I_filtered_10b[1566] = 046;
    I_filtered_10b[1565] = 035;
    I_filtered_10b[1564] = 021;
    I_filtered_10b[1563] = 00A;
    I_filtered_10b[1562] = 3F6;
    I_filtered_10b[1561] = 3E1;
    I_filtered_10b[1560] = 3CE;
    I_filtered_10b[1559] = 3C1;
    I_filtered_10b[1558] = 3B5;
    I_filtered_10b[1557] = 3AC;
    I_filtered_10b[1556] = 3A7;
    I_filtered_10b[1555] = 3A5;
    I_filtered_10b[1554] = 3A1;
    I_filtered_10b[1553] = 39F;
    I_filtered_10b[1552] = 39D;
    I_filtered_10b[1551] = 399;
    I_filtered_10b[1550] = 393;
    I_filtered_10b[1549] = 38C;
    I_filtered_10b[1548] = 381;
    I_filtered_10b[1547] = 378;
    I_filtered_10b[1546] = 36D;
    I_filtered_10b[1545] = 366;
    I_filtered_10b[1544] = 363;
    I_filtered_10b[1543] = 361;
    I_filtered_10b[1542] = 366;
    I_filtered_10b[1541] = 371;
    I_filtered_10b[1540] = 383;
    I_filtered_10b[1539] = 399;
    I_filtered_10b[1538] = 3B5;
    I_filtered_10b[1537] = 3D5;
    I_filtered_10b[1536] = 3F5;
    I_filtered_10b[1535] = 016;
    I_filtered_10b[1534] = 033;
    I_filtered_10b[1533] = 04B;
    I_filtered_10b[1532] = 05E;
    I_filtered_10b[1531] = 06B;
    I_filtered_10b[1530] = 071;
    I_filtered_10b[1529] = 06F;
    I_filtered_10b[1528] = 069;
    I_filtered_10b[1527] = 05D;
    I_filtered_10b[1526] = 04D;
    I_filtered_10b[1525] = 03B;
    I_filtered_10b[1524] = 026;
    I_filtered_10b[1523] = 013;
    I_filtered_10b[1522] = 003;
    I_filtered_10b[1521] = 3F6;
    I_filtered_10b[1520] = 3ED;
    I_filtered_10b[1519] = 3E5;
    I_filtered_10b[1518] = 3E1;
    I_filtered_10b[1517] = 3E0;
    I_filtered_10b[1516] = 3E1;
    I_filtered_10b[1515] = 3DF;
    I_filtered_10b[1514] = 3DC;
    I_filtered_10b[1513] = 3DB;
    I_filtered_10b[1512] = 3D4;
    I_filtered_10b[1511] = 3CD;
    I_filtered_10b[1510] = 3C3;
    I_filtered_10b[1509] = 3B8;
    I_filtered_10b[1508] = 3AE;
    I_filtered_10b[1507] = 3A5;
    I_filtered_10b[1506] = 39E;
    I_filtered_10b[1505] = 39C;
    I_filtered_10b[1504] = 39B;
    I_filtered_10b[1503] = 3A0;
    I_filtered_10b[1502] = 3A9;
    I_filtered_10b[1501] = 3B7;
    I_filtered_10b[1500] = 3C8;
    I_filtered_10b[1499] = 3DD;
    I_filtered_10b[1498] = 3F5;
    I_filtered_10b[1497] = 00B;
    I_filtered_10b[1496] = 022;
    I_filtered_10b[1495] = 036;
    I_filtered_10b[1494] = 045;
    I_filtered_10b[1493] = 052;
    I_filtered_10b[1492] = 05B;
    I_filtered_10b[1491] = 05F;
    I_filtered_10b[1490] = 05F;
    I_filtered_10b[1489] = 060;
    I_filtered_10b[1488] = 05D;
    I_filtered_10b[1487] = 05A;
    I_filtered_10b[1486] = 057;
    I_filtered_10b[1485] = 054;
    I_filtered_10b[1484] = 052;
    I_filtered_10b[1483] = 054;
    I_filtered_10b[1482] = 055;
    I_filtered_10b[1481] = 05A;
    I_filtered_10b[1480] = 05D;
    I_filtered_10b[1479] = 05E;
    I_filtered_10b[1478] = 05F;
    I_filtered_10b[1477] = 05E;
    I_filtered_10b[1476] = 056;
    I_filtered_10b[1475] = 049;
    I_filtered_10b[1474] = 03A;
    I_filtered_10b[1473] = 025;
    I_filtered_10b[1472] = 00C;
    I_filtered_10b[1471] = 3F1;
    I_filtered_10b[1470] = 3D4;
    I_filtered_10b[1469] = 3BA;
    I_filtered_10b[1468] = 3A6;
    I_filtered_10b[1467] = 395;
    I_filtered_10b[1466] = 38C;
    I_filtered_10b[1465] = 389;
    I_filtered_10b[1464] = 38F;
    I_filtered_10b[1463] = 39D;
    I_filtered_10b[1462] = 3B1;
    I_filtered_10b[1461] = 3CA;
    I_filtered_10b[1460] = 3E9;
    I_filtered_10b[1459] = 00A;
    I_filtered_10b[1458] = 02A;
    I_filtered_10b[1457] = 049;
    I_filtered_10b[1456] = 063;
    I_filtered_10b[1455] = 078;
    I_filtered_10b[1454] = 089;
    I_filtered_10b[1453] = 094;
    I_filtered_10b[1452] = 099;
    I_filtered_10b[1451] = 099;
    I_filtered_10b[1450] = 09A;
    I_filtered_10b[1449] = 097;
    I_filtered_10b[1448] = 091;
    I_filtered_10b[1447] = 08F;
    I_filtered_10b[1446] = 08C;
    I_filtered_10b[1445] = 08C;
    I_filtered_10b[1444] = 08E;
    I_filtered_10b[1443] = 090;
    I_filtered_10b[1442] = 093;
    I_filtered_10b[1441] = 095;
    I_filtered_10b[1440] = 093;
    I_filtered_10b[1439] = 093;
    I_filtered_10b[1438] = 08D;
    I_filtered_10b[1437] = 084;
    I_filtered_10b[1436] = 078;
    I_filtered_10b[1435] = 069;
    I_filtered_10b[1434] = 057;
    I_filtered_10b[1433] = 041;
    I_filtered_10b[1432] = 02D;
    I_filtered_10b[1431] = 017;
    I_filtered_10b[1430] = 004;
    I_filtered_10b[1429] = 3F7;
    I_filtered_10b[1428] = 3EB;
    I_filtered_10b[1427] = 3E1;
    I_filtered_10b[1426] = 3DA;
    I_filtered_10b[1425] = 3D9;
    I_filtered_10b[1424] = 3D5;
    I_filtered_10b[1423] = 3D3;
    I_filtered_10b[1422] = 3D1;
    I_filtered_10b[1421] = 3CE;
    I_filtered_10b[1420] = 3C8;
    I_filtered_10b[1419] = 3C0;
    I_filtered_10b[1418] = 3B6;
    I_filtered_10b[1417] = 3AB;
    I_filtered_10b[1416] = 3A1;
    I_filtered_10b[1415] = 399;
    I_filtered_10b[1414] = 396;
    I_filtered_10b[1413] = 395;
    I_filtered_10b[1412] = 39B;
    I_filtered_10b[1411] = 3A7;
    I_filtered_10b[1410] = 3BA;
    I_filtered_10b[1409] = 3CF;
    I_filtered_10b[1408] = 3EC;
    I_filtered_10b[1407] = 00C;
    I_filtered_10b[1406] = 02B;
    I_filtered_10b[1405] = 04B;
    I_filtered_10b[1404] = 067;
    I_filtered_10b[1403] = 07C;
    I_filtered_10b[1402] = 08E;
    I_filtered_10b[1401] = 09A;
    I_filtered_10b[1400] = 09F;
    I_filtered_10b[1399] = 09D;
    I_filtered_10b[1398] = 09A;
    I_filtered_10b[1397] = 092;
    I_filtered_10b[1396] = 088;
    I_filtered_10b[1395] = 07F;
    I_filtered_10b[1394] = 073;
    I_filtered_10b[1393] = 06A;
    I_filtered_10b[1392] = 066;
    I_filtered_10b[1391] = 061;
    I_filtered_10b[1390] = 062;
    I_filtered_10b[1389] = 061;
    I_filtered_10b[1388] = 05F;
    I_filtered_10b[1387] = 05F;
    I_filtered_10b[1386] = 05D;
    I_filtered_10b[1385] = 052;
    I_filtered_10b[1384] = 042;
    I_filtered_10b[1383] = 02F;
    I_filtered_10b[1382] = 013;
    I_filtered_10b[1381] = 3F6;
    I_filtered_10b[1380] = 3D4;
    I_filtered_10b[1379] = 3AE;
    I_filtered_10b[1378] = 38E;
    I_filtered_10b[1377] = 36F;
    I_filtered_10b[1376] = 358;
    I_filtered_10b[1375] = 34A;
    I_filtered_10b[1374] = 343;
    I_filtered_10b[1373] = 348;
    I_filtered_10b[1372] = 359;
    I_filtered_10b[1371] = 377;
    I_filtered_10b[1370] = 39C;
    I_filtered_10b[1369] = 3CB;
    I_filtered_10b[1368] = 3FE;
    I_filtered_10b[1367] = 031;
    I_filtered_10b[1366] = 067;
    I_filtered_10b[1365] = 094;
    I_filtered_10b[1364] = 0BD;
    I_filtered_10b[1363] = 0DB;
    I_filtered_10b[1362] = 0EF;
    I_filtered_10b[1361] = 0F6;
    I_filtered_10b[1360] = 0F4;
    I_filtered_10b[1359] = 0E6;
    I_filtered_10b[1358] = 0CB;
    I_filtered_10b[1357] = 0A7;
    I_filtered_10b[1356] = 07E;
    I_filtered_10b[1355] = 04F;
    I_filtered_10b[1354] = 020;
    I_filtered_10b[1353] = 3F2;
    I_filtered_10b[1352] = 3C8;
    I_filtered_10b[1351] = 3A5;
    I_filtered_10b[1350] = 38A;
    I_filtered_10b[1349] = 37A;
    I_filtered_10b[1348] = 377;
    I_filtered_10b[1347] = 37C;
    I_filtered_10b[1346] = 38D;
    I_filtered_10b[1345] = 3A8;
    I_filtered_10b[1344] = 3CB;
    I_filtered_10b[1343] = 3F4;
    I_filtered_10b[1342] = 021;
    I_filtered_10b[1341] = 04E;
    I_filtered_10b[1340] = 07A;
    I_filtered_10b[1339] = 0A2;
    I_filtered_10b[1338] = 0C4;
    I_filtered_10b[1337] = 0DE;
    I_filtered_10b[1336] = 0ED;
    I_filtered_10b[1335] = 0F0;
    I_filtered_10b[1334] = 0EC;
    I_filtered_10b[1333] = 0DC;
    I_filtered_10b[1332] = 0C2;
    I_filtered_10b[1331] = 09F;
    I_filtered_10b[1330] = 078;
    I_filtered_10b[1329] = 04B;
    I_filtered_10b[1328] = 01E;
    I_filtered_10b[1327] = 3F3;
    I_filtered_10b[1326] = 3CB;
    I_filtered_10b[1325] = 3AA;
    I_filtered_10b[1324] = 390;
    I_filtered_10b[1323] = 381;
    I_filtered_10b[1322] = 37D;
    I_filtered_10b[1321] = 382;
    I_filtered_10b[1320] = 390;
    I_filtered_10b[1319] = 3A6;
    I_filtered_10b[1318] = 3C4;
    I_filtered_10b[1317] = 3E5;
    I_filtered_10b[1316] = 00B;
    I_filtered_10b[1315] = 02F;
    I_filtered_10b[1314] = 051;
    I_filtered_10b[1313] = 070;
    I_filtered_10b[1312] = 087;
    I_filtered_10b[1311] = 09A;
    I_filtered_10b[1310] = 0A4;
    I_filtered_10b[1309] = 0A5;
    I_filtered_10b[1308] = 0A0;
    I_filtered_10b[1307] = 098;
    I_filtered_10b[1306] = 08C;
    I_filtered_10b[1305] = 07B;
    I_filtered_10b[1304] = 06C;
    I_filtered_10b[1303] = 05A;
    I_filtered_10b[1302] = 04D;
    I_filtered_10b[1301] = 041;
    I_filtered_10b[1300] = 036;
    I_filtered_10b[1299] = 02C;
    I_filtered_10b[1298] = 025;
    I_filtered_10b[1297] = 01D;
    I_filtered_10b[1296] = 01A;
    I_filtered_10b[1295] = 014;
    I_filtered_10b[1294] = 00D;
    I_filtered_10b[1293] = 006;
    I_filtered_10b[1292] = 3FF;
    I_filtered_10b[1291] = 3F5;
    I_filtered_10b[1290] = 3EC;
    I_filtered_10b[1289] = 3E4;
    I_filtered_10b[1288] = 3D8;
    I_filtered_10b[1287] = 3D0;
    I_filtered_10b[1286] = 3C5;
    I_filtered_10b[1285] = 3BE;
    I_filtered_10b[1284] = 3B5;
    I_filtered_10b[1283] = 3AD;
    I_filtered_10b[1282] = 3A6;
    I_filtered_10b[1281] = 39E;
    I_filtered_10b[1280] = 39B;
    I_filtered_10b[1279] = 397;
    I_filtered_10b[1278] = 394;
    I_filtered_10b[1277] = 390;
    I_filtered_10b[1276] = 38F;
    I_filtered_10b[1275] = 38D;
    I_filtered_10b[1274] = 38A;
    I_filtered_10b[1273] = 387;
    I_filtered_10b[1272] = 385;
    I_filtered_10b[1271] = 382;
    I_filtered_10b[1270] = 37F;
    I_filtered_10b[1269] = 37D;
    I_filtered_10b[1268] = 377;
    I_filtered_10b[1267] = 373;
    I_filtered_10b[1266] = 36D;
    I_filtered_10b[1265] = 366;
    I_filtered_10b[1264] = 35D;
    I_filtered_10b[1263] = 354;
    I_filtered_10b[1262] = 34B;
    I_filtered_10b[1261] = 342;
    I_filtered_10b[1260] = 33A;
    I_filtered_10b[1259] = 334;
    I_filtered_10b[1258] = 333;
    I_filtered_10b[1257] = 334;
    I_filtered_10b[1256] = 338;
    I_filtered_10b[1255] = 341;
    I_filtered_10b[1254] = 34E;
    I_filtered_10b[1253] = 35F;
    I_filtered_10b[1252] = 372;
    I_filtered_10b[1251] = 388;
    I_filtered_10b[1250] = 39C;
    I_filtered_10b[1249] = 3B2;
    I_filtered_10b[1248] = 3C6;
    I_filtered_10b[1247] = 3D7;
    I_filtered_10b[1246] = 3E5;
    I_filtered_10b[1245] = 3F1;
    I_filtered_10b[1244] = 3F8;
    I_filtered_10b[1243] = 3FC;
    I_filtered_10b[1242] = 3FD;
    I_filtered_10b[1241] = 3FA;
    I_filtered_10b[1240] = 3F6;
    I_filtered_10b[1239] = 3F0;
    I_filtered_10b[1238] = 3E9;
    I_filtered_10b[1237] = 3E0;
    I_filtered_10b[1236] = 3DC;
    I_filtered_10b[1235] = 3D7;
    I_filtered_10b[1234] = 3D8;
    I_filtered_10b[1233] = 3D7;
    I_filtered_10b[1232] = 3DB;
    I_filtered_10b[1231] = 3E0;
    I_filtered_10b[1230] = 3E7;
    I_filtered_10b[1229] = 3EE;
    I_filtered_10b[1228] = 3F2;
    I_filtered_10b[1227] = 3F9;
    I_filtered_10b[1226] = 3FC;
    I_filtered_10b[1225] = 000;
    I_filtered_10b[1224] = 000;
    I_filtered_10b[1223] = 000;
    I_filtered_10b[1222] = 001;
    I_filtered_10b[1221] = 003;
    I_filtered_10b[1220] = 004;
    I_filtered_10b[1219] = 009;
    I_filtered_10b[1218] = 00E;
    I_filtered_10b[1217] = 015;
    I_filtered_10b[1216] = 022;
    I_filtered_10b[1215] = 02E;
    I_filtered_10b[1214] = 03E;
    I_filtered_10b[1213] = 050;
    I_filtered_10b[1212] = 066;
    I_filtered_10b[1211] = 07A;
    I_filtered_10b[1210] = 08F;
    I_filtered_10b[1209] = 0A2;
    I_filtered_10b[1208] = 0B2;
    I_filtered_10b[1207] = 0BF;
    I_filtered_10b[1206] = 0C8;
    I_filtered_10b[1205] = 0CC;
    I_filtered_10b[1204] = 0CC;
    I_filtered_10b[1203] = 0CA;
    I_filtered_10b[1202] = 0C4;
    I_filtered_10b[1201] = 0BC;
    I_filtered_10b[1200] = 0B4;
    I_filtered_10b[1199] = 0AA;
    I_filtered_10b[1198] = 0A1;
    I_filtered_10b[1197] = 09B;
    I_filtered_10b[1196] = 095;
    I_filtered_10b[1195] = 094;
    I_filtered_10b[1194] = 092;
    I_filtered_10b[1193] = 08E;
    I_filtered_10b[1192] = 08D;
    I_filtered_10b[1191] = 08B;
    I_filtered_10b[1190] = 083;
    I_filtered_10b[1189] = 078;
    I_filtered_10b[1188] = 06A;
    I_filtered_10b[1187] = 057;
    I_filtered_10b[1186] = 040;
    I_filtered_10b[1185] = 027;
    I_filtered_10b[1184] = 00C;
    I_filtered_10b[1183] = 3F2;
    I_filtered_10b[1182] = 3DD;
    I_filtered_10b[1181] = 3CC;
    I_filtered_10b[1180] = 3C1;
    I_filtered_10b[1179] = 3BC;
    I_filtered_10b[1178] = 3C2;
    I_filtered_10b[1177] = 3CF;
    I_filtered_10b[1176] = 3E4;
    I_filtered_10b[1175] = 3FC;
    I_filtered_10b[1174] = 01C;
    I_filtered_10b[1173] = 03F;
    I_filtered_10b[1172] = 060;
    I_filtered_10b[1171] = 081;
    I_filtered_10b[1170] = 09C;
    I_filtered_10b[1169] = 0B2;
    I_filtered_10b[1168] = 0C4;
    I_filtered_10b[1167] = 0CF;
    I_filtered_10b[1166] = 0D2;
    I_filtered_10b[1165] = 0D2;
    I_filtered_10b[1164] = 0CF;
    I_filtered_10b[1163] = 0C8;
    I_filtered_10b[1162] = 0BD;
    I_filtered_10b[1161] = 0B5;
    I_filtered_10b[1160] = 0A9;
    I_filtered_10b[1159] = 0A0;
    I_filtered_10b[1158] = 09A;
    I_filtered_10b[1157] = 092;
    I_filtered_10b[1156] = 08F;
    I_filtered_10b[1155] = 08C;
    I_filtered_10b[1154] = 088;
    I_filtered_10b[1153] = 087;
    I_filtered_10b[1152] = 085;
    I_filtered_10b[1151] = 080;
    I_filtered_10b[1150] = 079;
    I_filtered_10b[1149] = 071;
    I_filtered_10b[1148] = 066;
    I_filtered_10b[1147] = 058;
    I_filtered_10b[1146] = 04A;
    I_filtered_10b[1145] = 039;
    I_filtered_10b[1144] = 02A;
    I_filtered_10b[1143] = 01E;
    I_filtered_10b[1142] = 014;
    I_filtered_10b[1141] = 00C;
    I_filtered_10b[1140] = 008;
    I_filtered_10b[1139] = 009;
    I_filtered_10b[1138] = 00C;
    I_filtered_10b[1137] = 013;
    I_filtered_10b[1136] = 01A;
    I_filtered_10b[1135] = 025;
    I_filtered_10b[1134] = 030;
    I_filtered_10b[1133] = 03B;
    I_filtered_10b[1132] = 043;
    I_filtered_10b[1131] = 04A;
    I_filtered_10b[1130] = 04C;
    I_filtered_10b[1129] = 04F;
    I_filtered_10b[1128] = 04F;
    I_filtered_10b[1127] = 04D;
    I_filtered_10b[1126] = 04B;
    I_filtered_10b[1125] = 04D;
    I_filtered_10b[1124] = 051;
    I_filtered_10b[1123] = 055;
    I_filtered_10b[1122] = 05E;
    I_filtered_10b[1121] = 067;
    I_filtered_10b[1120] = 074;
    I_filtered_10b[1119] = 082;
    I_filtered_10b[1118] = 08E;
    I_filtered_10b[1117] = 09A;
    I_filtered_10b[1116] = 0A3;
    I_filtered_10b[1115] = 0A5;
    I_filtered_10b[1114] = 0A5;
    I_filtered_10b[1113] = 09F;
    I_filtered_10b[1112] = 08F;
    I_filtered_10b[1111] = 079;
    I_filtered_10b[1110] = 05D;
    I_filtered_10b[1109] = 03A;
    I_filtered_10b[1108] = 011;
    I_filtered_10b[1107] = 3E8;
    I_filtered_10b[1106] = 3BD;
    I_filtered_10b[1105] = 396;
    I_filtered_10b[1104] = 377;
    I_filtered_10b[1103] = 35E;
    I_filtered_10b[1102] = 34F;
    I_filtered_10b[1101] = 349;
    I_filtered_10b[1100] = 350;
    I_filtered_10b[1099] = 35D;
    I_filtered_10b[1098] = 373;
    I_filtered_10b[1097] = 38F;
    I_filtered_10b[1096] = 3AF;
    I_filtered_10b[1095] = 3D1;
    I_filtered_10b[1094] = 3F0;
    I_filtered_10b[1093] = 00D;
    I_filtered_10b[1092] = 025;
    I_filtered_10b[1091] = 038;
    I_filtered_10b[1090] = 047;
    I_filtered_10b[1089] = 054;
    I_filtered_10b[1088] = 059;
    I_filtered_10b[1087] = 05E;
    I_filtered_10b[1086] = 066;
    I_filtered_10b[1085] = 06B;
    I_filtered_10b[1084] = 070;
    I_filtered_10b[1083] = 07A;
    I_filtered_10b[1082] = 085;
    I_filtered_10b[1081] = 090;
    I_filtered_10b[1080] = 0A0;
    I_filtered_10b[1079] = 0AC;
    I_filtered_10b[1078] = 0B8;
    I_filtered_10b[1077] = 0C2;
    I_filtered_10b[1076] = 0C8;
    I_filtered_10b[1075] = 0CC;
    I_filtered_10b[1074] = 0CB;
    I_filtered_10b[1073] = 0C7;
    I_filtered_10b[1072] = 0BD;
    I_filtered_10b[1071] = 0B2;
    I_filtered_10b[1070] = 0A4;
    I_filtered_10b[1069] = 096;
    I_filtered_10b[1068] = 08A;
    I_filtered_10b[1067] = 07B;
    I_filtered_10b[1066] = 071;
    I_filtered_10b[1065] = 066;
    I_filtered_10b[1064] = 05F;
    I_filtered_10b[1063] = 054;
    I_filtered_10b[1062] = 04D;
    I_filtered_10b[1061] = 045;
    I_filtered_10b[1060] = 03C;
    I_filtered_10b[1059] = 036;
    I_filtered_10b[1058] = 02E;
    I_filtered_10b[1057] = 027;
    I_filtered_10b[1056] = 01E;
    I_filtered_10b[1055] = 01A;
    I_filtered_10b[1054] = 011;
    I_filtered_10b[1053] = 00B;
    I_filtered_10b[1052] = 004;
    I_filtered_10b[1051] = 3FE;
    I_filtered_10b[1050] = 3F5;
    I_filtered_10b[1049] = 3EC;
    I_filtered_10b[1048] = 3E4;
    I_filtered_10b[1047] = 3D6;
    I_filtered_10b[1046] = 3CB;
    I_filtered_10b[1045] = 3BB;
    I_filtered_10b[1044] = 3AB;
    I_filtered_10b[1043] = 398;
    I_filtered_10b[1042] = 388;
    I_filtered_10b[1041] = 373;
    I_filtered_10b[1040] = 361;
    I_filtered_10b[1039] = 34E;
    I_filtered_10b[1038] = 340;
    I_filtered_10b[1037] = 335;
    I_filtered_10b[1036] = 32E;
    I_filtered_10b[1035] = 32B;
    I_filtered_10b[1034] = 32E;
    I_filtered_10b[1033] = 338;
    I_filtered_10b[1032] = 345;
    I_filtered_10b[1031] = 357;
    I_filtered_10b[1030] = 368;
    I_filtered_10b[1029] = 37B;
    I_filtered_10b[1028] = 390;
    I_filtered_10b[1027] = 3A1;
    I_filtered_10b[1026] = 3B1;
    I_filtered_10b[1025] = 3BD;
    I_filtered_10b[1024] = 3C7;
    I_filtered_10b[1023] = 3CB;
    I_filtered_10b[1022] = 3CD;
    I_filtered_10b[1021] = 3C7;
    I_filtered_10b[1020] = 3BB;
    I_filtered_10b[1019] = 3AD;
    I_filtered_10b[1018] = 398;
    I_filtered_10b[1017] = 383;
    I_filtered_10b[1016] = 369;
    I_filtered_10b[1015] = 350;
    I_filtered_10b[1014] = 33A;
    I_filtered_10b[1013] = 325;
    I_filtered_10b[1012] = 317;
    I_filtered_10b[1011] = 313;
    I_filtered_10b[1010] = 316;
    I_filtered_10b[1009] = 320;
    I_filtered_10b[1008] = 337;
    I_filtered_10b[1007] = 357;
    I_filtered_10b[1006] = 381;
    I_filtered_10b[1005] = 3B0;
    I_filtered_10b[1004] = 3E7;
    I_filtered_10b[1003] = 01C;
    I_filtered_10b[1002] = 055;
    I_filtered_10b[1001] = 088;
    I_filtered_10b[1000] = 0B6;
    I_filtered_10b[999] = 0D9;
    I_filtered_10b[998] = 0F1;
    I_filtered_10b[997] = 0FC;
    I_filtered_10b[996] = 0FB;
    I_filtered_10b[995] = 0EE;
    I_filtered_10b[994] = 0D2;
    I_filtered_10b[993] = 0AE;
    I_filtered_10b[992] = 082;
    I_filtered_10b[991] = 053;
    I_filtered_10b[990] = 022;
    I_filtered_10b[989] = 3F3;
    I_filtered_10b[988] = 3CB;
    I_filtered_10b[987] = 3A9;
    I_filtered_10b[986] = 38F;
    I_filtered_10b[985] = 380;
    I_filtered_10b[984] = 37D;
    I_filtered_10b[983] = 381;
    I_filtered_10b[982] = 38F;
    I_filtered_10b[981] = 3A5;
    I_filtered_10b[980] = 3C4;
    I_filtered_10b[979] = 3E5;
    I_filtered_10b[978] = 00C;
    I_filtered_10b[977] = 032;
    I_filtered_10b[976] = 056;
    I_filtered_10b[975] = 078;
    I_filtered_10b[974] = 092;
    I_filtered_10b[973] = 0A7;
    I_filtered_10b[972] = 0B1;
    I_filtered_10b[971] = 0B1;
    I_filtered_10b[970] = 0A9;
    I_filtered_10b[969] = 09A;
    I_filtered_10b[968] = 085;
    I_filtered_10b[967] = 069;
    I_filtered_10b[966] = 04C;
    I_filtered_10b[965] = 02A;
    I_filtered_10b[964] = 00D;
    I_filtered_10b[963] = 3F0;
    I_filtered_10b[962] = 3D6;
    I_filtered_10b[961] = 3C0;
    I_filtered_10b[960] = 3AE;
    I_filtered_10b[959] = 3A1;
    I_filtered_10b[958] = 39B;
    I_filtered_10b[957] = 397;
    I_filtered_10b[956] = 396;
    I_filtered_10b[955] = 399;
    I_filtered_10b[954] = 39F;
    I_filtered_10b[953] = 3A4;
    I_filtered_10b[952] = 3A9;
    I_filtered_10b[951] = 3AF;
    I_filtered_10b[950] = 3B3;
    I_filtered_10b[949] = 3B6;
    I_filtered_10b[948] = 3B9;
    I_filtered_10b[947] = 3BB;
    I_filtered_10b[946] = 3BB;
    I_filtered_10b[945] = 3B9;
    I_filtered_10b[944] = 3B8;
    I_filtered_10b[943] = 3B3;
    I_filtered_10b[942] = 3AE;
    I_filtered_10b[941] = 3A6;
    I_filtered_10b[940] = 39E;
    I_filtered_10b[939] = 395;
    I_filtered_10b[938] = 38B;
    I_filtered_10b[937] = 380;
    I_filtered_10b[936] = 376;
    I_filtered_10b[935] = 36B;
    I_filtered_10b[934] = 363;
    I_filtered_10b[933] = 361;
    I_filtered_10b[932] = 361;
    I_filtered_10b[931] = 365;
    I_filtered_10b[930] = 371;
    I_filtered_10b[929] = 383;
    I_filtered_10b[928] = 39A;
    I_filtered_10b[927] = 3B6;
    I_filtered_10b[926] = 3D6;
    I_filtered_10b[925] = 3F7;
    I_filtered_10b[924] = 01A;
    I_filtered_10b[923] = 03A;
    I_filtered_10b[922] = 055;
    I_filtered_10b[921] = 06A;
    I_filtered_10b[920] = 078;
    I_filtered_10b[919] = 07D;
    I_filtered_10b[918] = 079;
    I_filtered_10b[917] = 06D;
    I_filtered_10b[916] = 057;
    I_filtered_10b[915] = 03D;
    I_filtered_10b[914] = 01C;
    I_filtered_10b[913] = 3F9;
    I_filtered_10b[912] = 3D7;
    I_filtered_10b[911] = 3B4;
    I_filtered_10b[910] = 398;
    I_filtered_10b[909] = 37F;
    I_filtered_10b[908] = 36C;
    I_filtered_10b[907] = 35F;
    I_filtered_10b[906] = 35B;
    I_filtered_10b[905] = 35B;
    I_filtered_10b[904] = 361;
    I_filtered_10b[903] = 36D;
    I_filtered_10b[902] = 37E;
    I_filtered_10b[901] = 38F;
    I_filtered_10b[900] = 3A2;
    I_filtered_10b[899] = 3B5;
    I_filtered_10b[898] = 3C8;
    I_filtered_10b[897] = 3D9;
    I_filtered_10b[896] = 3E9;
    I_filtered_10b[895] = 3F4;
    I_filtered_10b[894] = 3FC;
    I_filtered_10b[893] = 3FE;
    I_filtered_10b[892] = 3FF;
    I_filtered_10b[891] = 3F9;
    I_filtered_10b[890] = 3EE;
    I_filtered_10b[889] = 3DF;
    I_filtered_10b[888] = 3CC;
    I_filtered_10b[887] = 3B5;
    I_filtered_10b[886] = 39B;
    I_filtered_10b[885] = 384;
    I_filtered_10b[884] = 36D;
    I_filtered_10b[883] = 35C;
    I_filtered_10b[882] = 34E;
    I_filtered_10b[881] = 34B;
    I_filtered_10b[880] = 34F;
    I_filtered_10b[879] = 35C;
    I_filtered_10b[878] = 373;
    I_filtered_10b[877] = 38F;
    I_filtered_10b[876] = 3B3;
    I_filtered_10b[875] = 3DA;
    I_filtered_10b[874] = 007;
    I_filtered_10b[873] = 02F;
    I_filtered_10b[872] = 05A;
    I_filtered_10b[871] = 07F;
    I_filtered_10b[870] = 09F;
    I_filtered_10b[869] = 0B9;
    I_filtered_10b[868] = 0CD;
    I_filtered_10b[867] = 0D8;
    I_filtered_10b[866] = 0DE;
    I_filtered_10b[865] = 0E1;
    I_filtered_10b[864] = 0DD;
    I_filtered_10b[863] = 0D6;
    I_filtered_10b[862] = 0CF;
    I_filtered_10b[861] = 0CA;
    I_filtered_10b[860] = 0C4;
    I_filtered_10b[859] = 0C0;
    I_filtered_10b[858] = 0BF;
    I_filtered_10b[857] = 0BD;
    I_filtered_10b[856] = 0BC;
    I_filtered_10b[855] = 0BA;
    I_filtered_10b[854] = 0BA;
    I_filtered_10b[853] = 0B6;
    I_filtered_10b[852] = 0B4;
    I_filtered_10b[851] = 0B1;
    I_filtered_10b[850] = 0AF;
    I_filtered_10b[849] = 0AC;
    I_filtered_10b[848] = 0A9;
    I_filtered_10b[847] = 0AA;
    I_filtered_10b[846] = 0A9;
    I_filtered_10b[845] = 0AA;
    I_filtered_10b[844] = 0AC;
    I_filtered_10b[843] = 0AD;
    I_filtered_10b[842] = 0A6;
    I_filtered_10b[841] = 09F;
    I_filtered_10b[840] = 094;
    I_filtered_10b[839] = 07F;
    I_filtered_10b[838] = 066;
    I_filtered_10b[837] = 046;
    I_filtered_10b[836] = 021;
    I_filtered_10b[835] = 3F4;
    I_filtered_10b[834] = 3C8;
    I_filtered_10b[833] = 399;
    I_filtered_10b[832] = 36D;
    I_filtered_10b[831] = 349;
    I_filtered_10b[830] = 32C;
    I_filtered_10b[829] = 319;
    I_filtered_10b[828] = 310;
    I_filtered_10b[827] = 315;
    I_filtered_10b[826] = 321;
    I_filtered_10b[825] = 337;
    I_filtered_10b[824] = 353;
    I_filtered_10b[823] = 374;
    I_filtered_10b[822] = 398;
    I_filtered_10b[821] = 3B8;
    I_filtered_10b[820] = 3D6;
    I_filtered_10b[819] = 3EE;
    I_filtered_10b[818] = 3FF;
    I_filtered_10b[817] = 00E;
    I_filtered_10b[816] = 01A;
    I_filtered_10b[815] = 020;
    I_filtered_10b[814] = 025;
    I_filtered_10b[813] = 02F;
    I_filtered_10b[812] = 039;
    I_filtered_10b[811] = 042;
    I_filtered_10b[810] = 053;
    I_filtered_10b[809] = 066;
    I_filtered_10b[808] = 07A;
    I_filtered_10b[807] = 092;
    I_filtered_10b[806] = 0A7;
    I_filtered_10b[805] = 0BA;
    I_filtered_10b[804] = 0C9;
    I_filtered_10b[803] = 0D2;
    I_filtered_10b[802] = 0D8;
    I_filtered_10b[801] = 0D5;
    I_filtered_10b[800] = 0CE;
    I_filtered_10b[799] = 0BF;
    I_filtered_10b[798] = 0AD;
    I_filtered_10b[797] = 096;
    I_filtered_10b[796] = 080;
    I_filtered_10b[795] = 06B;
    I_filtered_10b[794] = 054;
    I_filtered_10b[793] = 043;
    I_filtered_10b[792] = 034;
    I_filtered_10b[791] = 028;
    I_filtered_10b[790] = 01B;
    I_filtered_10b[789] = 014;
    I_filtered_10b[788] = 00B;
    I_filtered_10b[787] = 003;
    I_filtered_10b[786] = 3FD;
    I_filtered_10b[785] = 3F7;
    I_filtered_10b[784] = 3F0;
    I_filtered_10b[783] = 3E7;
    I_filtered_10b[782] = 3E2;
    I_filtered_10b[781] = 3D8;
    I_filtered_10b[780] = 3D1;
    I_filtered_10b[779] = 3C9;
    I_filtered_10b[778] = 3C3;
    I_filtered_10b[777] = 3BB;
    I_filtered_10b[776] = 3B3;
    I_filtered_10b[775] = 3AD;
    I_filtered_10b[774] = 3A3;
    I_filtered_10b[773] = 39B;
    I_filtered_10b[772] = 391;
    I_filtered_10b[771] = 386;
    I_filtered_10b[770] = 378;
    I_filtered_10b[769] = 36C;
    I_filtered_10b[768] = 35D;
    I_filtered_10b[767] = 34E;
    I_filtered_10b[766] = 340;
    I_filtered_10b[765] = 336;
    I_filtered_10b[764] = 330;
    I_filtered_10b[763] = 32E;
    I_filtered_10b[762] = 331;
    I_filtered_10b[761] = 339;
    I_filtered_10b[760] = 347;
    I_filtered_10b[759] = 358;
    I_filtered_10b[758] = 36D;
    I_filtered_10b[757] = 386;
    I_filtered_10b[756] = 39E;
    I_filtered_10b[755] = 3B6;
    I_filtered_10b[754] = 3CC;
    I_filtered_10b[753] = 3DC;
    I_filtered_10b[752] = 3E9;
    I_filtered_10b[751] = 3F4;
    I_filtered_10b[750] = 3F8;
    I_filtered_10b[749] = 3F8;
    I_filtered_10b[748] = 3F7;
    I_filtered_10b[747] = 3F4;
    I_filtered_10b[746] = 3F0;
    I_filtered_10b[745] = 3EC;
    I_filtered_10b[744] = 3E7;
    I_filtered_10b[743] = 3E4;
    I_filtered_10b[742] = 3E5;
    I_filtered_10b[741] = 3E6;
    I_filtered_10b[740] = 3EA;
    I_filtered_10b[739] = 3EC;
    I_filtered_10b[738] = 3EF;
    I_filtered_10b[737] = 3F2;
    I_filtered_10b[736] = 3F3;
    I_filtered_10b[735] = 3EE;
    I_filtered_10b[734] = 3E5;
    I_filtered_10b[733] = 3DB;
    I_filtered_10b[732] = 3CA;
    I_filtered_10b[731] = 3B9;
    I_filtered_10b[730] = 3A5;
    I_filtered_10b[729] = 38F;
    I_filtered_10b[728] = 37E;
    I_filtered_10b[727] = 36E;
    I_filtered_10b[726] = 362;
    I_filtered_10b[725] = 35C;
    I_filtered_10b[724] = 35B;
    I_filtered_10b[723] = 360;
    I_filtered_10b[722] = 36D;
    I_filtered_10b[721] = 380;
    I_filtered_10b[720] = 398;
    I_filtered_10b[719] = 3B4;
    I_filtered_10b[718] = 3D6;
    I_filtered_10b[717] = 3F7;
    I_filtered_10b[716] = 018;
    I_filtered_10b[715] = 036;
    I_filtered_10b[714] = 04D;
    I_filtered_10b[713] = 061;
    I_filtered_10b[712] = 06D;
    I_filtered_10b[711] = 071;
    I_filtered_10b[710] = 06E;
    I_filtered_10b[709] = 067;
    I_filtered_10b[708] = 05A;
    I_filtered_10b[707] = 04A;
    I_filtered_10b[706] = 039;
    I_filtered_10b[705] = 026;
    I_filtered_10b[704] = 016;
    I_filtered_10b[703] = 008;
    I_filtered_10b[702] = 3FD;
    I_filtered_10b[701] = 3F5;
    I_filtered_10b[700] = 3EE;
    I_filtered_10b[699] = 3E8;
    I_filtered_10b[698] = 3E6;
    I_filtered_10b[697] = 3E3;
    I_filtered_10b[696] = 3DD;
    I_filtered_10b[695] = 3D6;
    I_filtered_10b[694] = 3CF;
    I_filtered_10b[693] = 3C2;
    I_filtered_10b[692] = 3B6;
    I_filtered_10b[691] = 3A8;
    I_filtered_10b[690] = 397;
    I_filtered_10b[689] = 38A;
    I_filtered_10b[688] = 37D;
    I_filtered_10b[687] = 373;
    I_filtered_10b[686] = 36C;
    I_filtered_10b[685] = 367;
    I_filtered_10b[684] = 367;
    I_filtered_10b[683] = 36B;
    I_filtered_10b[682] = 375;
    I_filtered_10b[681] = 381;
    I_filtered_10b[680] = 391;
    I_filtered_10b[679] = 3A2;
    I_filtered_10b[678] = 3B4;
    I_filtered_10b[677] = 3C7;
    I_filtered_10b[676] = 3D6;
    I_filtered_10b[675] = 3E3;
    I_filtered_10b[674] = 3ED;
    I_filtered_10b[673] = 3F5;
    I_filtered_10b[672] = 3F8;
    I_filtered_10b[671] = 3F9;
    I_filtered_10b[670] = 3F5;
    I_filtered_10b[669] = 3EF;
    I_filtered_10b[668] = 3E6;
    I_filtered_10b[667] = 3DB;
    I_filtered_10b[666] = 3CF;
    I_filtered_10b[665] = 3C2;
    I_filtered_10b[664] = 3B7;
    I_filtered_10b[663] = 3AD;
    I_filtered_10b[662] = 3A6;
    I_filtered_10b[661] = 3A0;
    I_filtered_10b[660] = 39F;
    I_filtered_10b[659] = 3A1;
    I_filtered_10b[658] = 3A5;
    I_filtered_10b[657] = 3AD;
    I_filtered_10b[656] = 3B6;
    I_filtered_10b[655] = 3C3;
    I_filtered_10b[654] = 3D0;
    I_filtered_10b[653] = 3E1;
    I_filtered_10b[652] = 3EF;
    I_filtered_10b[651] = 3FD;
    I_filtered_10b[650] = 00B;
    I_filtered_10b[649] = 015;
    I_filtered_10b[648] = 01E;
    I_filtered_10b[647] = 023;
    I_filtered_10b[646] = 026;
    I_filtered_10b[645] = 024;
    I_filtered_10b[644] = 024;
    I_filtered_10b[643] = 022;
    I_filtered_10b[642] = 01F;
    I_filtered_10b[641] = 01E;
    I_filtered_10b[640] = 01C;
    I_filtered_10b[639] = 01D;
    I_filtered_10b[638] = 020;
    I_filtered_10b[637] = 023;
    I_filtered_10b[636] = 028;
    I_filtered_10b[635] = 02B;
    I_filtered_10b[634] = 02B;
    I_filtered_10b[633] = 02C;
    I_filtered_10b[632] = 028;
    I_filtered_10b[631] = 01F;
    I_filtered_10b[630] = 012;
    I_filtered_10b[629] = 002;
    I_filtered_10b[628] = 3ED;
    I_filtered_10b[627] = 3D4;
    I_filtered_10b[626] = 3B9;
    I_filtered_10b[625] = 39F;
    I_filtered_10b[624] = 386;
    I_filtered_10b[623] = 374;
    I_filtered_10b[622] = 365;
    I_filtered_10b[621] = 35D;
    I_filtered_10b[620] = 35B;
    I_filtered_10b[619] = 362;
    I_filtered_10b[618] = 36C;
    I_filtered_10b[617] = 37C;
    I_filtered_10b[616] = 38F;
    I_filtered_10b[615] = 3A5;
    I_filtered_10b[614] = 3BD;
    I_filtered_10b[613] = 3D1;
    I_filtered_10b[612] = 3E5;
    I_filtered_10b[611] = 3F5;
    I_filtered_10b[610] = 000;
    I_filtered_10b[609] = 00B;
    I_filtered_10b[608] = 014;
    I_filtered_10b[607] = 01A;
    I_filtered_10b[606] = 01F;
    I_filtered_10b[605] = 029;
    I_filtered_10b[604] = 034;
    I_filtered_10b[603] = 040;
    I_filtered_10b[602] = 051;
    I_filtered_10b[601] = 064;
    I_filtered_10b[600] = 077;
    I_filtered_10b[599] = 091;
    I_filtered_10b[598] = 0A5;
    I_filtered_10b[597] = 0BC;
    I_filtered_10b[596] = 0CC;
    I_filtered_10b[595] = 0D7;
    I_filtered_10b[594] = 0DE;
    I_filtered_10b[593] = 0DE;
    I_filtered_10b[592] = 0D5;
    I_filtered_10b[591] = 0C2;
    I_filtered_10b[590] = 0AA;
    I_filtered_10b[589] = 08A;
    I_filtered_10b[588] = 069;
    I_filtered_10b[587] = 045;
    I_filtered_10b[586] = 01F;
    I_filtered_10b[585] = 000;
    I_filtered_10b[584] = 3E2;
    I_filtered_10b[583] = 3CC;
    I_filtered_10b[582] = 3BD;
    I_filtered_10b[581] = 3B6;
    I_filtered_10b[580] = 3B7;
    I_filtered_10b[579] = 3C2;
    I_filtered_10b[578] = 3D8;
    I_filtered_10b[577] = 3F4;
    I_filtered_10b[576] = 017;
    I_filtered_10b[575] = 03D;
    I_filtered_10b[574] = 067;
    I_filtered_10b[573] = 090;
    I_filtered_10b[572] = 0B4;
    I_filtered_10b[571] = 0D4;
    I_filtered_10b[570] = 0EB;
    I_filtered_10b[569] = 0F6;
    I_filtered_10b[568] = 0F6;
    I_filtered_10b[567] = 0ED;
    I_filtered_10b[566] = 0D6;
    I_filtered_10b[565] = 0B4;
    I_filtered_10b[564] = 087;
    I_filtered_10b[563] = 055;
    I_filtered_10b[562] = 019;
    I_filtered_10b[561] = 3E0;
    I_filtered_10b[560] = 3A6;
    I_filtered_10b[559] = 370;
    I_filtered_10b[558] = 344;
    I_filtered_10b[557] = 321;
    I_filtered_10b[556] = 30B;
    I_filtered_10b[555] = 304;
    I_filtered_10b[554] = 309;
    I_filtered_10b[553] = 319;
    I_filtered_10b[552] = 335;
    I_filtered_10b[551] = 359;
    I_filtered_10b[550] = 383;
    I_filtered_10b[549] = 3B2;
    I_filtered_10b[548] = 3DE;
    I_filtered_10b[547] = 007;
    I_filtered_10b[546] = 02C;
    I_filtered_10b[545] = 048;
    I_filtered_10b[544] = 05F;
    I_filtered_10b[543] = 06E;
    I_filtered_10b[542] = 071;
    I_filtered_10b[541] = 070;
    I_filtered_10b[540] = 06B;
    I_filtered_10b[539] = 062;
    I_filtered_10b[538] = 054;
    I_filtered_10b[537] = 049;
    I_filtered_10b[536] = 03D;
    I_filtered_10b[535] = 033;
    I_filtered_10b[534] = 02C;
    I_filtered_10b[533] = 026;
    I_filtered_10b[532] = 020;
    I_filtered_10b[531] = 01D;
    I_filtered_10b[530] = 019;
    I_filtered_10b[529] = 01A;
    I_filtered_10b[528] = 017;
    I_filtered_10b[527] = 014;
    I_filtered_10b[526] = 011;
    I_filtered_10b[525] = 00F;
    I_filtered_10b[524] = 009;
    I_filtered_10b[523] = 004;
    I_filtered_10b[522] = 000;
    I_filtered_10b[521] = 3FB;
    I_filtered_10b[520] = 3F8;
    I_filtered_10b[519] = 3F6;
    I_filtered_10b[518] = 3F4;
    I_filtered_10b[517] = 3F0;
    I_filtered_10b[516] = 3EC;
    I_filtered_10b[515] = 3E9;
    I_filtered_10b[514] = 3E1;
    I_filtered_10b[513] = 3D9;
    I_filtered_10b[512] = 3CE;
    I_filtered_10b[511] = 3C2;
    I_filtered_10b[510] = 3B4;
    I_filtered_10b[509] = 3A6;
    I_filtered_10b[508] = 395;
    I_filtered_10b[507] = 386;
    I_filtered_10b[506] = 377;
    I_filtered_10b[505] = 36C;
    I_filtered_10b[504] = 365;
    I_filtered_10b[503] = 361;
    I_filtered_10b[502] = 362;
    I_filtered_10b[501] = 36A;
    I_filtered_10b[500] = 378;
    I_filtered_10b[499] = 38A;
    I_filtered_10b[498] = 3A1;
    I_filtered_10b[497] = 3BA;
    I_filtered_10b[496] = 3D4;
    I_filtered_10b[495] = 3F0;
    I_filtered_10b[494] = 007;
    I_filtered_10b[493] = 01D;
    I_filtered_10b[492] = 02D;
    I_filtered_10b[491] = 039;
    I_filtered_10b[490] = 03E;
    I_filtered_10b[489] = 03D;
    I_filtered_10b[488] = 035;
    I_filtered_10b[487] = 024;
    I_filtered_10b[486] = 010;
    I_filtered_10b[485] = 3F6;
    I_filtered_10b[484] = 3D7;
    I_filtered_10b[483] = 3B5;
    I_filtered_10b[482] = 397;
    I_filtered_10b[481] = 37A;
    I_filtered_10b[480] = 365;
    I_filtered_10b[479] = 353;
    I_filtered_10b[478] = 34D;
    I_filtered_10b[477] = 34F;
    I_filtered_10b[476] = 35A;
    I_filtered_10b[475] = 36D;
    I_filtered_10b[474] = 386;
    I_filtered_10b[473] = 3A6;
    I_filtered_10b[472] = 3C8;
    I_filtered_10b[471] = 3EF;
    I_filtered_10b[470] = 00F;
    I_filtered_10b[469] = 032;
    I_filtered_10b[468] = 050;
    I_filtered_10b[467] = 06A;
    I_filtered_10b[466] = 07F;
    I_filtered_10b[465] = 090;
    I_filtered_10b[464] = 099;
    I_filtered_10b[463] = 09F;
    I_filtered_10b[462] = 0A5;
    I_filtered_10b[461] = 0A5;
    I_filtered_10b[460] = 0A4;
    I_filtered_10b[459] = 0A5;
    I_filtered_10b[458] = 0A6;
    I_filtered_10b[457] = 0A6;
    I_filtered_10b[456] = 0AB;
    I_filtered_10b[455] = 0AE;
    I_filtered_10b[454] = 0B4;
    I_filtered_10b[453] = 0B8;
    I_filtered_10b[452] = 0BC;
    I_filtered_10b[451] = 0C0;
    I_filtered_10b[450] = 0C2;
    I_filtered_10b[449] = 0C2;
    I_filtered_10b[448] = 0BE;
    I_filtered_10b[447] = 0BA;
    I_filtered_10b[446] = 0B3;
    I_filtered_10b[445] = 0AE;
    I_filtered_10b[444] = 0A7;
    I_filtered_10b[443] = 09E;
    I_filtered_10b[442] = 099;
    I_filtered_10b[441] = 092;
    I_filtered_10b[440] = 08E;
    I_filtered_10b[439] = 086;
    I_filtered_10b[438] = 081;
    I_filtered_10b[437] = 07B;
    I_filtered_10b[436] = 076;
    I_filtered_10b[435] = 074;
    I_filtered_10b[434] = 070;
    I_filtered_10b[433] = 06F;
    I_filtered_10b[432] = 06B;
    I_filtered_10b[431] = 06C;
    I_filtered_10b[430] = 06C;
    I_filtered_10b[429] = 06A;
    I_filtered_10b[428] = 06B;
    I_filtered_10b[427] = 06A;
    I_filtered_10b[426] = 065;
    I_filtered_10b[425] = 05F;
    I_filtered_10b[424] = 059;
    I_filtered_10b[423] = 04C;
    I_filtered_10b[422] = 03B;
    I_filtered_10b[421] = 026;
    I_filtered_10b[420] = 00D;
    I_filtered_10b[419] = 3EF;
    I_filtered_10b[418] = 3D0;
    I_filtered_10b[417] = 3AE;
    I_filtered_10b[416] = 38D;
    I_filtered_10b[415] = 372;
    I_filtered_10b[414] = 35C;
    I_filtered_10b[413] = 34F;
    I_filtered_10b[412] = 349;
    I_filtered_10b[411] = 34F;
    I_filtered_10b[410] = 35F;
    I_filtered_10b[409] = 378;
    I_filtered_10b[408] = 397;
    I_filtered_10b[407] = 3BE;
    I_filtered_10b[406] = 3EA;
    I_filtered_10b[405] = 014;
    I_filtered_10b[404] = 03D;
    I_filtered_10b[403] = 061;
    I_filtered_10b[402] = 07C;
    I_filtered_10b[401] = 092;
    I_filtered_10b[400] = 0A0;
    I_filtered_10b[399] = 0A5;
    I_filtered_10b[398] = 0A2;
    I_filtered_10b[397] = 09E;
    I_filtered_10b[396] = 096;
    I_filtered_10b[395] = 089;
    I_filtered_10b[394] = 07F;
    I_filtered_10b[393] = 073;
    I_filtered_10b[392] = 06C;
    I_filtered_10b[391] = 068;
    I_filtered_10b[390] = 064;
    I_filtered_10b[389] = 064;
    I_filtered_10b[388] = 063;
    I_filtered_10b[387] = 060;
    I_filtered_10b[386] = 05F;
    I_filtered_10b[385] = 05A;
    I_filtered_10b[384] = 04F;
    I_filtered_10b[383] = 03E;
    I_filtered_10b[382] = 02C;
    I_filtered_10b[381] = 011;
    I_filtered_10b[380] = 3F6;
    I_filtered_10b[379] = 3DA;
    I_filtered_10b[378] = 3B8;
    I_filtered_10b[377] = 39D;
    I_filtered_10b[376] = 382;
    I_filtered_10b[375] = 36E;
    I_filtered_10b[374] = 35E;
    I_filtered_10b[373] = 355;
    I_filtered_10b[372] = 353;
    I_filtered_10b[371] = 359;
    I_filtered_10b[370] = 36A;
    I_filtered_10b[369] = 37E;
    I_filtered_10b[368] = 399;
    I_filtered_10b[367] = 3B5;
    I_filtered_10b[366] = 3D5;
    I_filtered_10b[365] = 3F4;
    I_filtered_10b[364] = 00E;
    I_filtered_10b[363] = 025;
    I_filtered_10b[362] = 037;
    I_filtered_10b[361] = 041;
    I_filtered_10b[360] = 044;
    I_filtered_10b[359] = 041;
    I_filtered_10b[358] = 034;
    I_filtered_10b[357] = 01F;
    I_filtered_10b[356] = 004;
    I_filtered_10b[355] = 3E4;
    I_filtered_10b[354] = 3C0;
    I_filtered_10b[353] = 39A;
    I_filtered_10b[352] = 374;
    I_filtered_10b[351] = 353;
    I_filtered_10b[350] = 334;
    I_filtered_10b[349] = 31E;
    I_filtered_10b[348] = 312;
    I_filtered_10b[347] = 310;
    I_filtered_10b[346] = 316;
    I_filtered_10b[345] = 329;
    I_filtered_10b[344] = 346;
    I_filtered_10b[343] = 36D;
    I_filtered_10b[342] = 399;
    I_filtered_10b[341] = 3CE;
    I_filtered_10b[340] = 002;
    I_filtered_10b[339] = 036;
    I_filtered_10b[338] = 067;
    I_filtered_10b[337] = 08D;
    I_filtered_10b[336] = 0AC;
    I_filtered_10b[335] = 0BE;
    I_filtered_10b[334] = 0C3;
    I_filtered_10b[333] = 0BB;
    I_filtered_10b[332] = 0AA;
    I_filtered_10b[331] = 08E;
    I_filtered_10b[330] = 06B;
    I_filtered_10b[329] = 043;
    I_filtered_10b[328] = 017;
    I_filtered_10b[327] = 3EF;
    I_filtered_10b[326] = 3C8;
    I_filtered_10b[325] = 3A7;
    I_filtered_10b[324] = 38C;
    I_filtered_10b[323] = 376;
    I_filtered_10b[322] = 367;
    I_filtered_10b[321] = 361;
    I_filtered_10b[320] = 35E;
    I_filtered_10b[319] = 35D;
    I_filtered_10b[318] = 361;
    I_filtered_10b[317] = 369;
    I_filtered_10b[316] = 36E;
    I_filtered_10b[315] = 373;
    I_filtered_10b[314] = 378;
    I_filtered_10b[313] = 37A;
    I_filtered_10b[312] = 37D;
    I_filtered_10b[311] = 37F;
    I_filtered_10b[310] = 380;
    I_filtered_10b[309] = 381;
    I_filtered_10b[308] = 37F;
    I_filtered_10b[307] = 380;
    I_filtered_10b[306] = 37E;
    I_filtered_10b[305] = 37D;
    I_filtered_10b[304] = 37A;
    I_filtered_10b[303] = 378;
    I_filtered_10b[302] = 376;
    I_filtered_10b[301] = 372;
    I_filtered_10b[300] = 36E;
    I_filtered_10b[299] = 36A;
    I_filtered_10b[298] = 365;
    I_filtered_10b[297] = 362;
    I_filtered_10b[296] = 364;
    I_filtered_10b[295] = 367;
    I_filtered_10b[294] = 36D;
    I_filtered_10b[293] = 37A;
    I_filtered_10b[292] = 38B;
    I_filtered_10b[291] = 3A1;
    I_filtered_10b[290] = 3BA;
    I_filtered_10b[289] = 3D7;
    I_filtered_10b[288] = 3F2;
    I_filtered_10b[287] = 012;
    I_filtered_10b[286] = 02E;
    I_filtered_10b[285] = 04A;
    I_filtered_10b[284] = 05E;
    I_filtered_10b[283] = 06E;
    I_filtered_10b[282] = 077;
    I_filtered_10b[281] = 079;
    I_filtered_10b[280] = 073;
    I_filtered_10b[279] = 062;
    I_filtered_10b[278] = 04D;
    I_filtered_10b[277] = 031;
    I_filtered_10b[276] = 013;
    I_filtered_10b[275] = 3F1;
    I_filtered_10b[274] = 3D1;
    I_filtered_10b[273] = 3B5;
    I_filtered_10b[272] = 39D;
    I_filtered_10b[271] = 38B;
    I_filtered_10b[270] = 383;
    I_filtered_10b[269] = 383;
    I_filtered_10b[268] = 38A;
    I_filtered_10b[267] = 39B;
    I_filtered_10b[266] = 3B4;
    I_filtered_10b[265] = 3D5;
    I_filtered_10b[264] = 3FA;
    I_filtered_10b[263] = 023;
    I_filtered_10b[262] = 04B;
    I_filtered_10b[261] = 075;
    I_filtered_10b[260] = 099;
    I_filtered_10b[259] = 0BB;
    I_filtered_10b[258] = 0D4;
    I_filtered_10b[257] = 0E4;
    I_filtered_10b[256] = 0EA;
    I_filtered_10b[255] = 0E9;
    I_filtered_10b[254] = 0DE;
    I_filtered_10b[253] = 0C9;
    I_filtered_10b[252] = 0AC;
    I_filtered_10b[251] = 08B;
    I_filtered_10b[250] = 066;
    I_filtered_10b[249] = 040;
    I_filtered_10b[248] = 01B;
    I_filtered_10b[247] = 3FA;
    I_filtered_10b[246] = 3DD;
    I_filtered_10b[245] = 3C7;
    I_filtered_10b[244] = 3BA;
    I_filtered_10b[243] = 3B6;
    I_filtered_10b[242] = 3BA;
    I_filtered_10b[241] = 3C7;
    I_filtered_10b[240] = 3DD;
    I_filtered_10b[239] = 3FA;
    I_filtered_10b[238] = 01B;
    I_filtered_10b[237] = 041;
    I_filtered_10b[236] = 068;
    I_filtered_10b[235] = 08D;
    I_filtered_10b[234] = 0AF;
    I_filtered_10b[233] = 0CB;
    I_filtered_10b[232] = 0E0;
    I_filtered_10b[231] = 0EA;
    I_filtered_10b[230] = 0EA;
    I_filtered_10b[229] = 0E2;
    I_filtered_10b[228] = 0D1;
    I_filtered_10b[227] = 0B8;
    I_filtered_10b[226] = 096;
    I_filtered_10b[225] = 073;
    I_filtered_10b[224] = 04A;
    I_filtered_10b[223] = 025;
    I_filtered_10b[222] = 3FF;
    I_filtered_10b[221] = 3DD;
    I_filtered_10b[220] = 3BF;
    I_filtered_10b[219] = 3A8;
    I_filtered_10b[218] = 397;
    I_filtered_10b[217] = 38F;
    I_filtered_10b[216] = 38C;
    I_filtered_10b[215] = 38D;
    I_filtered_10b[214] = 396;
    I_filtered_10b[213] = 3A3;
    I_filtered_10b[212] = 3B1;
    I_filtered_10b[211] = 3BF;
    I_filtered_10b[210] = 3CF;
    I_filtered_10b[209] = 3DC;
    I_filtered_10b[208] = 3E8;
    I_filtered_10b[207] = 3F1;
    I_filtered_10b[206] = 3F8;
    I_filtered_10b[205] = 3FB;
    I_filtered_10b[204] = 3F8;
    I_filtered_10b[203] = 3F6;
    I_filtered_10b[202] = 3ED;
    I_filtered_10b[201] = 3E3;
    I_filtered_10b[200] = 3D5;
    I_filtered_10b[199] = 3C6;
    I_filtered_10b[198] = 3B5;
    I_filtered_10b[197] = 3A4;
    I_filtered_10b[196] = 391;
    I_filtered_10b[195] = 381;
    I_filtered_10b[194] = 36F;
    I_filtered_10b[193] = 363;
    I_filtered_10b[192] = 35D;
    I_filtered_10b[191] = 35B;
    I_filtered_10b[190] = 35E;
    I_filtered_10b[189] = 369;
    I_filtered_10b[188] = 37C;
    I_filtered_10b[187] = 395;
    I_filtered_10b[186] = 3B2;
    I_filtered_10b[185] = 3D6;
    I_filtered_10b[184] = 3FC;
    I_filtered_10b[183] = 020;
    I_filtered_10b[182] = 044;
    I_filtered_10b[181] = 05F;
    I_filtered_10b[180] = 075;
    I_filtered_10b[179] = 081;
    I_filtered_10b[178] = 083;
    I_filtered_10b[177] = 07A;
    I_filtered_10b[176] = 068;
    I_filtered_10b[175] = 04E;
    I_filtered_10b[174] = 02E;
    I_filtered_10b[173] = 008;
    I_filtered_10b[172] = 3DF;
    I_filtered_10b[171] = 3BA;
    I_filtered_10b[170] = 394;
    I_filtered_10b[169] = 375;
    I_filtered_10b[168] = 35A;
    I_filtered_10b[167] = 345;
    I_filtered_10b[166] = 335;
    I_filtered_10b[165] = 32E;
    I_filtered_10b[164] = 329;
    I_filtered_10b[163] = 327;
    I_filtered_10b[162] = 32A;
    I_filtered_10b[161] = 331;
    I_filtered_10b[160] = 336;
    I_filtered_10b[159] = 33A;
    I_filtered_10b[158] = 33E;
    I_filtered_10b[157] = 341;
    I_filtered_10b[156] = 344;
    I_filtered_10b[155] = 347;
    I_filtered_10b[154] = 349;
    I_filtered_10b[153] = 34C;
    I_filtered_10b[152] = 34C;
    I_filtered_10b[151] = 34F;
    I_filtered_10b[150] = 34E;
    I_filtered_10b[149] = 34C;
    I_filtered_10b[148] = 34A;
    I_filtered_10b[147] = 345;
    I_filtered_10b[146] = 33F;
    I_filtered_10b[145] = 334;
    I_filtered_10b[144] = 32C;
    I_filtered_10b[143] = 322;
    I_filtered_10b[142] = 31A;
    I_filtered_10b[141] = 315;
    I_filtered_10b[140] = 31A;
    I_filtered_10b[139] = 322;
    I_filtered_10b[138] = 331;
    I_filtered_10b[137] = 34A;
    I_filtered_10b[136] = 368;
    I_filtered_10b[135] = 38F;
    I_filtered_10b[134] = 3B9;
    I_filtered_10b[133] = 3EB;
    I_filtered_10b[132] = 016;
    I_filtered_10b[131] = 048;
    I_filtered_10b[130] = 074;
    I_filtered_10b[129] = 09C;
    I_filtered_10b[128] = 0BB;
    I_filtered_10b[127] = 0D5;
    I_filtered_10b[126] = 0E4;
    I_filtered_10b[125] = 0EB;
    I_filtered_10b[124] = 0ED;
    I_filtered_10b[123] = 0E3;
    I_filtered_10b[122] = 0D7;
    I_filtered_10b[121] = 0C5;
    I_filtered_10b[120] = 0B6;
    I_filtered_10b[119] = 0A3;
    I_filtered_10b[118] = 093;
    I_filtered_10b[117] = 088;
    I_filtered_10b[116] = 07E;
    I_filtered_10b[115] = 078;
    I_filtered_10b[114] = 073;
    I_filtered_10b[113] = 075;
    I_filtered_10b[112] = 075;
    I_filtered_10b[111] = 07A;
    I_filtered_10b[110] = 081;
    I_filtered_10b[109] = 08B;
    I_filtered_10b[108] = 095;
    I_filtered_10b[107] = 0A2;
    I_filtered_10b[106] = 0B0;
    I_filtered_10b[105] = 0BE;
    I_filtered_10b[104] = 0CB;
    I_filtered_10b[103] = 0D9;
    I_filtered_10b[102] = 0E2;
    I_filtered_10b[101] = 0E2;
    I_filtered_10b[100] = 0DE;
    I_filtered_10b[99] = 0D5;
    I_filtered_10b[98] = 0C1;
    I_filtered_10b[97] = 0A7;
    I_filtered_10b[96] = 084;
    I_filtered_10b[95] = 05D;
    I_filtered_10b[94] = 02E;
    I_filtered_10b[93] = 001;
    I_filtered_10b[92] = 3D1;
    I_filtered_10b[91] = 3A5;
    I_filtered_10b[90] = 37F;
    I_filtered_10b[89] = 361;
    I_filtered_10b[88] = 34D;
    I_filtered_10b[87] = 343;
    I_filtered_10b[86] = 346;
    I_filtered_10b[85] = 351;
    I_filtered_10b[84] = 368;
    I_filtered_10b[83] = 385;
    I_filtered_10b[82] = 3A8;
    I_filtered_10b[81] = 3CE;
    I_filtered_10b[80] = 3F4;
    I_filtered_10b[79] = 016;
    I_filtered_10b[78] = 034;
    I_filtered_10b[77] = 04B;
    I_filtered_10b[76] = 05D;
    I_filtered_10b[75] = 069;
    I_filtered_10b[74] = 06B;
    I_filtered_10b[73] = 06A;
    I_filtered_10b[72] = 066;
    I_filtered_10b[71] = 05E;
    I_filtered_10b[70] = 052;
    I_filtered_10b[69] = 048;
    I_filtered_10b[68] = 03C;
    I_filtered_10b[67] = 033;
    I_filtered_10b[66] = 02B;
    I_filtered_10b[65] = 023;
    I_filtered_10b[64] = 01C;
    I_filtered_10b[63] = 018;
    I_filtered_10b[62] = 014;
    I_filtered_10b[61] = 014;
    I_filtered_10b[60] = 012;
    I_filtered_10b[59] = 012;
    I_filtered_10b[58] = 013;
    I_filtered_10b[57] = 016;
    I_filtered_10b[56] = 018;
    I_filtered_10b[55] = 01C;
    I_filtered_10b[54] = 020;
    I_filtered_10b[53] = 024;
    I_filtered_10b[52] = 029;
    I_filtered_10b[51] = 02D;
    I_filtered_10b[50] = 030;
    I_filtered_10b[49] = 02F;
    I_filtered_10b[48] = 02C;
    I_filtered_10b[47] = 026;
    I_filtered_10b[46] = 01B;
    I_filtered_10b[45] = 00E;
    I_filtered_10b[44] = 3FD;
    I_filtered_10b[43] = 3EA;
    I_filtered_10b[42] = 3D2;
    I_filtered_10b[41] = 3BC;
    I_filtered_10b[40] = 3A3;
    I_filtered_10b[39] = 38D;
    I_filtered_10b[38] = 37A;
    I_filtered_10b[37] = 36C;
    I_filtered_10b[36] = 362;
    I_filtered_10b[35] = 35E;
    I_filtered_10b[34] = 360;
    I_filtered_10b[33] = 368;
    I_filtered_10b[32] = 375;
    I_filtered_10b[31] = 385;
    I_filtered_10b[30] = 399;
    I_filtered_10b[29] = 3AF;
    I_filtered_10b[28] = 3C4;
    I_filtered_10b[27] = 3D9;
    I_filtered_10b[26] = 3EA;
    I_filtered_10b[25] = 3F8;
    I_filtered_10b[24] = 003;
    I_filtered_10b[23] = 00C;
    I_filtered_10b[22] = 00F;
    I_filtered_10b[21] = 010;
    I_filtered_10b[20] = 010;
    I_filtered_10b[19] = 00D;
    I_filtered_10b[18] = 009;
    I_filtered_10b[17] = 006;
    I_filtered_10b[16] = 002;
    I_filtered_10b[15] = 3FF;
    I_filtered_10b[14] = 3FE;
    I_filtered_10b[13] = 3FC;
    I_filtered_10b[12] = 3FC;
    I_filtered_10b[11] = 3FC;
    I_filtered_10b[10] = 3FE;
    I_filtered_10b[9] = 000;
    I_filtered_10b[8] = 001;
    I_filtered_10b[7] = 002;
    I_filtered_10b[6] = 002;
    I_filtered_10b[5] = 004;
    I_filtered_10b[4] = 002;
    I_filtered_10b[3] = 002;
    I_filtered_10b[2] = 001;
    I_filtered_10b[1] = 000;
    I_filtered_10b[0] = 000;


// Q Channel 10b Expected output
    Q_filtered_10b[1733] = 000;
    Q_filtered_10b[1732] = 000;
    Q_filtered_10b[1731] = 000;
    Q_filtered_10b[1730] = 000;
    Q_filtered_10b[1729] = 000;
    Q_filtered_10b[1728] = 000;
    Q_filtered_10b[1727] = 000;
    Q_filtered_10b[1726] = 000;
    Q_filtered_10b[1725] = 000;
    Q_filtered_10b[1724] = 000;
    Q_filtered_10b[1723] = 000;
    Q_filtered_10b[1722] = 000;
    Q_filtered_10b[1721] = 000;
    Q_filtered_10b[1720] = 000;
    Q_filtered_10b[1719] = 001;
    Q_filtered_10b[1718] = 002;
    Q_filtered_10b[1717] = 002;
    Q_filtered_10b[1716] = 004;
    Q_filtered_10b[1715] = 002;
    Q_filtered_10b[1714] = 002;
    Q_filtered_10b[1713] = 001;
    Q_filtered_10b[1712] = 000;
    Q_filtered_10b[1711] = 3FE;
    Q_filtered_10b[1710] = 3FC;
    Q_filtered_10b[1709] = 3FC;
    Q_filtered_10b[1708] = 3FC;
    Q_filtered_10b[1707] = 3FE;
    Q_filtered_10b[1706] = 3FE;
    Q_filtered_10b[1705] = 001;
    Q_filtered_10b[1704] = 005;
    Q_filtered_10b[1703] = 006;
    Q_filtered_10b[1702] = 00B;
    Q_filtered_10b[1701] = 00D;
    Q_filtered_10b[1700] = 00E;
    Q_filtered_10b[1699] = 00E;
    Q_filtered_10b[1698] = 00B;
    Q_filtered_10b[1697] = 005;
    Q_filtered_10b[1696] = 3FB;
    Q_filtered_10b[1695] = 3EE;
    Q_filtered_10b[1694] = 3DD;
    Q_filtered_10b[1693] = 3CA;
    Q_filtered_10b[1692] = 3B4;
    Q_filtered_10b[1691] = 39F;
    Q_filtered_10b[1690] = 38C;
    Q_filtered_10b[1689] = 37C;
    Q_filtered_10b[1688] = 36F;
    Q_filtered_10b[1687] = 369;
    Q_filtered_10b[1686] = 369;
    Q_filtered_10b[1685] = 36F;
    Q_filtered_10b[1684] = 37D;
    Q_filtered_10b[1683] = 38E;
    Q_filtered_10b[1682] = 3A4;
    Q_filtered_10b[1681] = 3BD;
    Q_filtered_10b[1680] = 3D8;
    Q_filtered_10b[1679] = 3F1;
    Q_filtered_10b[1678] = 00A;
    Q_filtered_10b[1677] = 020;
    Q_filtered_10b[1676] = 033;
    Q_filtered_10b[1675] = 041;
    Q_filtered_10b[1674] = 04E;
    Q_filtered_10b[1673] = 055;
    Q_filtered_10b[1672] = 05C;
    Q_filtered_10b[1671] = 060;
    Q_filtered_10b[1670] = 061;
    Q_filtered_10b[1669] = 061;
    Q_filtered_10b[1668] = 064;
    Q_filtered_10b[1667] = 066;
    Q_filtered_10b[1666] = 067;
    Q_filtered_10b[1665] = 06B;
    Q_filtered_10b[1664] = 06F;
    Q_filtered_10b[1663] = 071;
    Q_filtered_10b[1662] = 074;
    Q_filtered_10b[1661] = 077;
    Q_filtered_10b[1660] = 078;
    Q_filtered_10b[1659] = 079;
    Q_filtered_10b[1658] = 079;
    Q_filtered_10b[1657] = 079;
    Q_filtered_10b[1656] = 07A;
    Q_filtered_10b[1655] = 07C;
    Q_filtered_10b[1654] = 07D;
    Q_filtered_10b[1653] = 081;
    Q_filtered_10b[1652] = 086;
    Q_filtered_10b[1651] = 088;
    Q_filtered_10b[1650] = 08F;
    Q_filtered_10b[1649] = 093;
    Q_filtered_10b[1648] = 093;
    Q_filtered_10b[1647] = 08E;
    Q_filtered_10b[1646] = 089;
    Q_filtered_10b[1645] = 07A;
    Q_filtered_10b[1644] = 067;
    Q_filtered_10b[1643] = 04F;
    Q_filtered_10b[1642] = 031;
    Q_filtered_10b[1641] = 011;
    Q_filtered_10b[1640] = 3F0;
    Q_filtered_10b[1639] = 3CB;
    Q_filtered_10b[1638] = 3AC;
    Q_filtered_10b[1637] = 38D;
    Q_filtered_10b[1636] = 376;
    Q_filtered_10b[1635] = 364;
    Q_filtered_10b[1634] = 35C;
    Q_filtered_10b[1633] = 359;
    Q_filtered_10b[1632] = 362;
    Q_filtered_10b[1631] = 376;
    Q_filtered_10b[1630] = 38F;
    Q_filtered_10b[1629] = 3AE;
    Q_filtered_10b[1628] = 3D1;
    Q_filtered_10b[1627] = 3F9;
    Q_filtered_10b[1626] = 01D;
    Q_filtered_10b[1625] = 03C;
    Q_filtered_10b[1624] = 057;
    Q_filtered_10b[1623] = 06B;
    Q_filtered_10b[1622] = 076;
    Q_filtered_10b[1621] = 076;
    Q_filtered_10b[1620] = 071;
    Q_filtered_10b[1619] = 061;
    Q_filtered_10b[1618] = 04A;
    Q_filtered_10b[1617] = 02A;
    Q_filtered_10b[1616] = 008;
    Q_filtered_10b[1615] = 3E0;
    Q_filtered_10b[1614] = 3B7;
    Q_filtered_10b[1613] = 392;
    Q_filtered_10b[1612] = 36F;
    Q_filtered_10b[1611] = 352;
    Q_filtered_10b[1610] = 33C;
    Q_filtered_10b[1609] = 32F;
    Q_filtered_10b[1608] = 32E;
    Q_filtered_10b[1607] = 331;
    Q_filtered_10b[1606] = 33F;
    Q_filtered_10b[1605] = 352;
    Q_filtered_10b[1604] = 36D;
    Q_filtered_10b[1603] = 387;
    Q_filtered_10b[1602] = 3A8;
    Q_filtered_10b[1601] = 3C8;
    Q_filtered_10b[1600] = 3E3;
    Q_filtered_10b[1599] = 3FF;
    Q_filtered_10b[1598] = 011;
    Q_filtered_10b[1597] = 021;
    Q_filtered_10b[1596] = 02A;
    Q_filtered_10b[1595] = 02D;
    Q_filtered_10b[1594] = 02B;
    Q_filtered_10b[1593] = 028;
    Q_filtered_10b[1592] = 025;
    Q_filtered_10b[1591] = 01E;
    Q_filtered_10b[1590] = 01D;
    Q_filtered_10b[1589] = 01A;
    Q_filtered_10b[1588] = 01B;
    Q_filtered_10b[1587] = 01F;
    Q_filtered_10b[1586] = 021;
    Q_filtered_10b[1585] = 027;
    Q_filtered_10b[1584] = 02A;
    Q_filtered_10b[1583] = 02C;
    Q_filtered_10b[1582] = 02D;
    Q_filtered_10b[1581] = 028;
    Q_filtered_10b[1580] = 01E;
    Q_filtered_10b[1579] = 00E;
    Q_filtered_10b[1578] = 3FC;
    Q_filtered_10b[1577] = 3E1;
    Q_filtered_10b[1576] = 3C6;
    Q_filtered_10b[1575] = 3A7;
    Q_filtered_10b[1574] = 389;
    Q_filtered_10b[1573] = 36F;
    Q_filtered_10b[1572] = 359;
    Q_filtered_10b[1571] = 348;
    Q_filtered_10b[1570] = 33C;
    Q_filtered_10b[1569] = 339;
    Q_filtered_10b[1568] = 33A;
    Q_filtered_10b[1567] = 343;
    Q_filtered_10b[1566] = 351;
    Q_filtered_10b[1565] = 364;
    Q_filtered_10b[1564] = 378;
    Q_filtered_10b[1563] = 390;
    Q_filtered_10b[1562] = 3A7;
    Q_filtered_10b[1561] = 3BC;
    Q_filtered_10b[1560] = 3D0;
    Q_filtered_10b[1559] = 3DD;
    Q_filtered_10b[1558] = 3E8;
    Q_filtered_10b[1557] = 3F0;
    Q_filtered_10b[1556] = 3F4;
    Q_filtered_10b[1555] = 3F5;
    Q_filtered_10b[1554] = 3F7;
    Q_filtered_10b[1553] = 3F8;
    Q_filtered_10b[1552] = 3F8;
    Q_filtered_10b[1551] = 3FC;
    Q_filtered_10b[1550] = 3FD;
    Q_filtered_10b[1549] = 001;
    Q_filtered_10b[1548] = 009;
    Q_filtered_10b[1547] = 00E;
    Q_filtered_10b[1546] = 017;
    Q_filtered_10b[1545] = 01C;
    Q_filtered_10b[1544] = 022;
    Q_filtered_10b[1543] = 027;
    Q_filtered_10b[1542] = 029;
    Q_filtered_10b[1541] = 026;
    Q_filtered_10b[1540] = 01E;
    Q_filtered_10b[1539] = 014;
    Q_filtered_10b[1538] = 004;
    Q_filtered_10b[1537] = 3F4;
    Q_filtered_10b[1536] = 3DF;
    Q_filtered_10b[1535] = 3CA;
    Q_filtered_10b[1534] = 3BB;
    Q_filtered_10b[1533] = 3AB;
    Q_filtered_10b[1532] = 3A0;
    Q_filtered_10b[1531] = 39A;
    Q_filtered_10b[1530] = 39A;
    Q_filtered_10b[1529] = 39E;
    Q_filtered_10b[1528] = 3AA;
    Q_filtered_10b[1527] = 3BB;
    Q_filtered_10b[1526] = 3D2;
    Q_filtered_10b[1525] = 3EC;
    Q_filtered_10b[1524] = 009;
    Q_filtered_10b[1523] = 027;
    Q_filtered_10b[1522] = 045;
    Q_filtered_10b[1521] = 05E;
    Q_filtered_10b[1520] = 077;
    Q_filtered_10b[1519] = 088;
    Q_filtered_10b[1518] = 095;
    Q_filtered_10b[1517] = 099;
    Q_filtered_10b[1516] = 09A;
    Q_filtered_10b[1515] = 092;
    Q_filtered_10b[1514] = 084;
    Q_filtered_10b[1513] = 070;
    Q_filtered_10b[1512] = 05A;
    Q_filtered_10b[1511] = 03F;
    Q_filtered_10b[1510] = 021;
    Q_filtered_10b[1509] = 008;
    Q_filtered_10b[1508] = 3F0;
    Q_filtered_10b[1507] = 3DE;
    Q_filtered_10b[1506] = 3CF;
    Q_filtered_10b[1505] = 3C8;
    Q_filtered_10b[1504] = 3C8;
    Q_filtered_10b[1503] = 3CE;
    Q_filtered_10b[1502] = 3D9;
    Q_filtered_10b[1501] = 3E8;
    Q_filtered_10b[1500] = 3FC;
    Q_filtered_10b[1499] = 010;
    Q_filtered_10b[1498] = 027;
    Q_filtered_10b[1497] = 03D;
    Q_filtered_10b[1496] = 050;
    Q_filtered_10b[1495] = 062;
    Q_filtered_10b[1494] = 070;
    Q_filtered_10b[1493] = 07A;
    Q_filtered_10b[1492] = 082;
    Q_filtered_10b[1491] = 083;
    Q_filtered_10b[1490] = 085;
    Q_filtered_10b[1489] = 084;
    Q_filtered_10b[1488] = 083;
    Q_filtered_10b[1487] = 07E;
    Q_filtered_10b[1486] = 07F;
    Q_filtered_10b[1485] = 07D;
    Q_filtered_10b[1484] = 07D;
    Q_filtered_10b[1483] = 07E;
    Q_filtered_10b[1482] = 07E;
    Q_filtered_10b[1481] = 07F;
    Q_filtered_10b[1480] = 080;
    Q_filtered_10b[1479] = 080;
    Q_filtered_10b[1478] = 07E;
    Q_filtered_10b[1477] = 07C;
    Q_filtered_10b[1476] = 076;
    Q_filtered_10b[1475] = 06F;
    Q_filtered_10b[1474] = 067;
    Q_filtered_10b[1473] = 05C;
    Q_filtered_10b[1472] = 051;
    Q_filtered_10b[1471] = 046;
    Q_filtered_10b[1470] = 03A;
    Q_filtered_10b[1469] = 02E;
    Q_filtered_10b[1468] = 026;
    Q_filtered_10b[1467] = 01E;
    Q_filtered_10b[1466] = 017;
    Q_filtered_10b[1465] = 011;
    Q_filtered_10b[1464] = 00E;
    Q_filtered_10b[1463] = 00A;
    Q_filtered_10b[1462] = 009;
    Q_filtered_10b[1461] = 006;
    Q_filtered_10b[1460] = 003;
    Q_filtered_10b[1459] = 000;
    Q_filtered_10b[1458] = 3FD;
    Q_filtered_10b[1457] = 3F8;
    Q_filtered_10b[1456] = 3F3;
    Q_filtered_10b[1455] = 3EC;
    Q_filtered_10b[1454] = 3E7;
    Q_filtered_10b[1453] = 3E2;
    Q_filtered_10b[1452] = 3DE;
    Q_filtered_10b[1451] = 3DC;
    Q_filtered_10b[1450] = 3DD;
    Q_filtered_10b[1449] = 3E2;
    Q_filtered_10b[1448] = 3E7;
    Q_filtered_10b[1447] = 3F0;
    Q_filtered_10b[1446] = 3F8;
    Q_filtered_10b[1445] = 003;
    Q_filtered_10b[1444] = 00E;
    Q_filtered_10b[1443] = 015;
    Q_filtered_10b[1442] = 01E;
    Q_filtered_10b[1441] = 023;
    Q_filtered_10b[1440] = 027;
    Q_filtered_10b[1439] = 027;
    Q_filtered_10b[1438] = 026;
    Q_filtered_10b[1437] = 021;
    Q_filtered_10b[1436] = 018;
    Q_filtered_10b[1435] = 00D;
    Q_filtered_10b[1434] = 3FF;
    Q_filtered_10b[1433] = 3ED;
    Q_filtered_10b[1432] = 3DA;
    Q_filtered_10b[1431] = 3C9;
    Q_filtered_10b[1430] = 3B8;
    Q_filtered_10b[1429] = 3AC;
    Q_filtered_10b[1428] = 3A2;
    Q_filtered_10b[1427] = 39E;
    Q_filtered_10b[1426] = 3A0;
    Q_filtered_10b[1425] = 3A6;
    Q_filtered_10b[1424] = 3B1;
    Q_filtered_10b[1423] = 3BE;
    Q_filtered_10b[1422] = 3D0;
    Q_filtered_10b[1421] = 3E2;
    Q_filtered_10b[1420] = 3F5;
    Q_filtered_10b[1419] = 005;
    Q_filtered_10b[1418] = 015;
    Q_filtered_10b[1417] = 024;
    Q_filtered_10b[1416] = 031;
    Q_filtered_10b[1415] = 03A;
    Q_filtered_10b[1414] = 044;
    Q_filtered_10b[1413] = 04A;
    Q_filtered_10b[1412] = 053;
    Q_filtered_10b[1411] = 05A;
    Q_filtered_10b[1410] = 060;
    Q_filtered_10b[1409] = 066;
    Q_filtered_10b[1408] = 070;
    Q_filtered_10b[1407] = 07B;
    Q_filtered_10b[1406] = 084;
    Q_filtered_10b[1405] = 08E;
    Q_filtered_10b[1404] = 098;
    Q_filtered_10b[1403] = 09F;
    Q_filtered_10b[1402] = 0A5;
    Q_filtered_10b[1401] = 0AA;
    Q_filtered_10b[1400] = 0AC;
    Q_filtered_10b[1399] = 0AD;
    Q_filtered_10b[1398] = 0AC;
    Q_filtered_10b[1397] = 0AC;
    Q_filtered_10b[1396] = 0AC;
    Q_filtered_10b[1395] = 0AE;
    Q_filtered_10b[1394] = 0B0;
    Q_filtered_10b[1393] = 0B5;
    Q_filtered_10b[1392] = 0BB;
    Q_filtered_10b[1391] = 0BE;
    Q_filtered_10b[1390] = 0C5;
    Q_filtered_10b[1389] = 0C9;
    Q_filtered_10b[1388] = 0C8;
    Q_filtered_10b[1387] = 0C2;
    Q_filtered_10b[1386] = 0B9;
    Q_filtered_10b[1385] = 0A6;
    Q_filtered_10b[1384] = 090;
    Q_filtered_10b[1383] = 073;
    Q_filtered_10b[1382] = 051;
    Q_filtered_10b[1381] = 02C;
    Q_filtered_10b[1380] = 008;
    Q_filtered_10b[1379] = 3E0;
    Q_filtered_10b[1378] = 3BD;
    Q_filtered_10b[1377] = 39B;
    Q_filtered_10b[1376] = 383;
    Q_filtered_10b[1375] = 36D;
    Q_filtered_10b[1374] = 361;
    Q_filtered_10b[1373] = 35B;
    Q_filtered_10b[1372] = 35D;
    Q_filtered_10b[1371] = 36A;
    Q_filtered_10b[1370] = 37A;
    Q_filtered_10b[1369] = 38E;
    Q_filtered_10b[1368] = 3A5;
    Q_filtered_10b[1367] = 3C1;
    Q_filtered_10b[1366] = 3D7;
    Q_filtered_10b[1365] = 3EA;
    Q_filtered_10b[1364] = 3F8;
    Q_filtered_10b[1363] = 003;
    Q_filtered_10b[1362] = 007;
    Q_filtered_10b[1361] = 004;
    Q_filtered_10b[1360] = 3FE;
    Q_filtered_10b[1359] = 3F2;
    Q_filtered_10b[1358] = 3E4;
    Q_filtered_10b[1357] = 3D0;
    Q_filtered_10b[1356] = 3BC;
    Q_filtered_10b[1355] = 3A4;
    Q_filtered_10b[1354] = 38D;
    Q_filtered_10b[1353] = 379;
    Q_filtered_10b[1352] = 365;
    Q_filtered_10b[1351] = 355;
    Q_filtered_10b[1350] = 349;
    Q_filtered_10b[1349] = 342;
    Q_filtered_10b[1348] = 344;
    Q_filtered_10b[1347] = 346;
    Q_filtered_10b[1346] = 34E;
    Q_filtered_10b[1345] = 357;
    Q_filtered_10b[1344] = 365;
    Q_filtered_10b[1343] = 370;
    Q_filtered_10b[1342] = 37D;
    Q_filtered_10b[1341] = 387;
    Q_filtered_10b[1340] = 391;
    Q_filtered_10b[1339] = 39B;
    Q_filtered_10b[1338] = 3A2;
    Q_filtered_10b[1337] = 3A8;
    Q_filtered_10b[1336] = 3AF;
    Q_filtered_10b[1335] = 3B6;
    Q_filtered_10b[1334] = 3BC;
    Q_filtered_10b[1333] = 3C6;
    Q_filtered_10b[1332] = 3CF;
    Q_filtered_10b[1331] = 3DB;
    Q_filtered_10b[1330] = 3EA;
    Q_filtered_10b[1329] = 3F8;
    Q_filtered_10b[1328] = 005;
    Q_filtered_10b[1327] = 016;
    Q_filtered_10b[1326] = 025;
    Q_filtered_10b[1325] = 035;
    Q_filtered_10b[1324] = 040;
    Q_filtered_10b[1323] = 04C;
    Q_filtered_10b[1322] = 055;
    Q_filtered_10b[1321] = 05D;
    Q_filtered_10b[1320] = 060;
    Q_filtered_10b[1319] = 05E;
    Q_filtered_10b[1318] = 05C;
    Q_filtered_10b[1317] = 057;
    Q_filtered_10b[1316] = 053;
    Q_filtered_10b[1315] = 04A;
    Q_filtered_10b[1314] = 043;
    Q_filtered_10b[1313] = 03F;
    Q_filtered_10b[1312] = 03B;
    Q_filtered_10b[1311] = 038;
    Q_filtered_10b[1310] = 038;
    Q_filtered_10b[1309] = 03A;
    Q_filtered_10b[1308] = 03E;
    Q_filtered_10b[1307] = 044;
    Q_filtered_10b[1306] = 04D;
    Q_filtered_10b[1305] = 059;
    Q_filtered_10b[1304] = 067;
    Q_filtered_10b[1303] = 078;
    Q_filtered_10b[1302] = 08B;
    Q_filtered_10b[1301] = 09C;
    Q_filtered_10b[1300] = 0AC;
    Q_filtered_10b[1299] = 0B8;
    Q_filtered_10b[1298] = 0C2;
    Q_filtered_10b[1297] = 0C6;
    Q_filtered_10b[1296] = 0C2;
    Q_filtered_10b[1295] = 0BA;
    Q_filtered_10b[1294] = 0AC;
    Q_filtered_10b[1293] = 09C;
    Q_filtered_10b[1292] = 086;
    Q_filtered_10b[1291] = 070;
    Q_filtered_10b[1290] = 055;
    Q_filtered_10b[1289] = 03E;
    Q_filtered_10b[1288] = 028;
    Q_filtered_10b[1287] = 011;
    Q_filtered_10b[1286] = 003;
    Q_filtered_10b[1285] = 3F7;
    Q_filtered_10b[1284] = 3EB;
    Q_filtered_10b[1283] = 3E4;
    Q_filtered_10b[1282] = 3DF;
    Q_filtered_10b[1281] = 3D6;
    Q_filtered_10b[1280] = 3CE;
    Q_filtered_10b[1279] = 3C4;
    Q_filtered_10b[1278] = 3B3;
    Q_filtered_10b[1277] = 3A4;
    Q_filtered_10b[1276] = 391;
    Q_filtered_10b[1275] = 379;
    Q_filtered_10b[1274] = 366;
    Q_filtered_10b[1273] = 34E;
    Q_filtered_10b[1272] = 33E;
    Q_filtered_10b[1271] = 332;
    Q_filtered_10b[1270] = 32E;
    Q_filtered_10b[1269] = 32F;
    Q_filtered_10b[1268] = 33E;
    Q_filtered_10b[1267] = 357;
    Q_filtered_10b[1266] = 376;
    Q_filtered_10b[1265] = 3A0;
    Q_filtered_10b[1264] = 3CA;
    Q_filtered_10b[1263] = 3FA;
    Q_filtered_10b[1262] = 02B;
    Q_filtered_10b[1261] = 052;
    Q_filtered_10b[1260] = 078;
    Q_filtered_10b[1259] = 094;
    Q_filtered_10b[1258] = 0A8;
    Q_filtered_10b[1257] = 0AF;
    Q_filtered_10b[1256] = 0B0;
    Q_filtered_10b[1255] = 0A3;
    Q_filtered_10b[1254] = 08A;
    Q_filtered_10b[1253] = 06A;
    Q_filtered_10b[1252] = 044;
    Q_filtered_10b[1251] = 01A;
    Q_filtered_10b[1250] = 3EB;
    Q_filtered_10b[1249] = 3BF;
    Q_filtered_10b[1248] = 39B;
    Q_filtered_10b[1247] = 379;
    Q_filtered_10b[1246] = 360;
    Q_filtered_10b[1245] = 352;
    Q_filtered_10b[1244] = 351;
    Q_filtered_10b[1243] = 355;
    Q_filtered_10b[1242] = 368;
    Q_filtered_10b[1241] = 383;
    Q_filtered_10b[1240] = 3A9;
    Q_filtered_10b[1239] = 3D2;
    Q_filtered_10b[1238] = 004;
    Q_filtered_10b[1237] = 039;
    Q_filtered_10b[1236] = 068;
    Q_filtered_10b[1235] = 094;
    Q_filtered_10b[1234] = 0B8;
    Q_filtered_10b[1233] = 0D4;
    Q_filtered_10b[1232] = 0E3;
    Q_filtered_10b[1231] = 0E3;
    Q_filtered_10b[1230] = 0DA;
    Q_filtered_10b[1229] = 0C5;
    Q_filtered_10b[1228] = 0A9;
    Q_filtered_10b[1227] = 082;
    Q_filtered_10b[1226] = 05C;
    Q_filtered_10b[1225] = 02F;
    Q_filtered_10b[1224] = 005;
    Q_filtered_10b[1223] = 3DF;
    Q_filtered_10b[1222] = 3BB;
    Q_filtered_10b[1221] = 39F;
    Q_filtered_10b[1220] = 38A;
    Q_filtered_10b[1219] = 378;
    Q_filtered_10b[1218] = 372;
    Q_filtered_10b[1217] = 36C;
    Q_filtered_10b[1216] = 369;
    Q_filtered_10b[1215] = 36A;
    Q_filtered_10b[1214] = 36E;
    Q_filtered_10b[1213] = 36A;
    Q_filtered_10b[1212] = 36A;
    Q_filtered_10b[1211] = 368;
    Q_filtered_10b[1210] = 362;
    Q_filtered_10b[1209] = 35E;
    Q_filtered_10b[1208] = 358;
    Q_filtered_10b[1207] = 354;
    Q_filtered_10b[1206] = 350;
    Q_filtered_10b[1205] = 34F;
    Q_filtered_10b[1204] = 34F;
    Q_filtered_10b[1203] = 354;
    Q_filtered_10b[1202] = 35B;
    Q_filtered_10b[1201] = 363;
    Q_filtered_10b[1200] = 36F;
    Q_filtered_10b[1199] = 37A;
    Q_filtered_10b[1198] = 385;
    Q_filtered_10b[1197] = 391;
    Q_filtered_10b[1196] = 39B;
    Q_filtered_10b[1195] = 3A1;
    Q_filtered_10b[1194] = 3A7;
    Q_filtered_10b[1193] = 3AE;
    Q_filtered_10b[1192] = 3B6;
    Q_filtered_10b[1191] = 3BB;
    Q_filtered_10b[1190] = 3C5;
    Q_filtered_10b[1189] = 3CE;
    Q_filtered_10b[1188] = 3DB;
    Q_filtered_10b[1187] = 3EA;
    Q_filtered_10b[1186] = 3FB;
    Q_filtered_10b[1185] = 00D;
    Q_filtered_10b[1184] = 020;
    Q_filtered_10b[1183] = 033;
    Q_filtered_10b[1182] = 044;
    Q_filtered_10b[1181] = 051;
    Q_filtered_10b[1180] = 05B;
    Q_filtered_10b[1179] = 060;
    Q_filtered_10b[1178] = 060;
    Q_filtered_10b[1177] = 05B;
    Q_filtered_10b[1176] = 051;
    Q_filtered_10b[1175] = 045;
    Q_filtered_10b[1174] = 035;
    Q_filtered_10b[1173] = 024;
    Q_filtered_10b[1172] = 012;
    Q_filtered_10b[1171] = 003;
    Q_filtered_10b[1170] = 3F6;
    Q_filtered_10b[1169] = 3EF;
    Q_filtered_10b[1168] = 3E8;
    Q_filtered_10b[1167] = 3E4;
    Q_filtered_10b[1166] = 3E4;
    Q_filtered_10b[1165] = 3E4;
    Q_filtered_10b[1164] = 3E3;
    Q_filtered_10b[1163] = 3E1;
    Q_filtered_10b[1162] = 3DF;
    Q_filtered_10b[1161] = 3D8;
    Q_filtered_10b[1160] = 3D2;
    Q_filtered_10b[1159] = 3C7;
    Q_filtered_10b[1158] = 3BC;
    Q_filtered_10b[1157] = 3B3;
    Q_filtered_10b[1156] = 3A9;
    Q_filtered_10b[1155] = 3A2;
    Q_filtered_10b[1154] = 39F;
    Q_filtered_10b[1153] = 3A0;
    Q_filtered_10b[1152] = 3A5;
    Q_filtered_10b[1151] = 3B1;
    Q_filtered_10b[1150] = 3C1;
    Q_filtered_10b[1149] = 3D5;
    Q_filtered_10b[1148] = 3EF;
    Q_filtered_10b[1147] = 00B;
    Q_filtered_10b[1146] = 028;
    Q_filtered_10b[1145] = 044;
    Q_filtered_10b[1144] = 05D;
    Q_filtered_10b[1143] = 070;
    Q_filtered_10b[1142] = 080;
    Q_filtered_10b[1141] = 08B;
    Q_filtered_10b[1140] = 08E;
    Q_filtered_10b[1139] = 08E;
    Q_filtered_10b[1138] = 08A;
    Q_filtered_10b[1137] = 083;
    Q_filtered_10b[1136] = 07A;
    Q_filtered_10b[1135] = 073;
    Q_filtered_10b[1134] = 068;
    Q_filtered_10b[1133] = 060;
    Q_filtered_10b[1132] = 05C;
    Q_filtered_10b[1131] = 056;
    Q_filtered_10b[1130] = 058;
    Q_filtered_10b[1129] = 057;
    Q_filtered_10b[1128] = 056;
    Q_filtered_10b[1127] = 055;
    Q_filtered_10b[1126] = 054;
    Q_filtered_10b[1125] = 04A;
    Q_filtered_10b[1124] = 03C;
    Q_filtered_10b[1123] = 02B;
    Q_filtered_10b[1122] = 011;
    Q_filtered_10b[1121] = 3F8;
    Q_filtered_10b[1120] = 3DA;
    Q_filtered_10b[1119] = 3B8;
    Q_filtered_10b[1118] = 39D;
    Q_filtered_10b[1117] = 380;
    Q_filtered_10b[1116] = 36B;
    Q_filtered_10b[1115] = 35C;
    Q_filtered_10b[1114] = 356;
    Q_filtered_10b[1113] = 357;
    Q_filtered_10b[1112] = 366;
    Q_filtered_10b[1111] = 381;
    Q_filtered_10b[1110] = 3A2;
    Q_filtered_10b[1109] = 3CE;
    Q_filtered_10b[1108] = 3FB;
    Q_filtered_10b[1107] = 02F;
    Q_filtered_10b[1106] = 062;
    Q_filtered_10b[1105] = 08C;
    Q_filtered_10b[1104] = 0B4;
    Q_filtered_10b[1103] = 0D1;
    Q_filtered_10b[1102] = 0E4;
    Q_filtered_10b[1101] = 0E8;
    Q_filtered_10b[1100] = 0E5;
    Q_filtered_10b[1099] = 0D1;
    Q_filtered_10b[1098] = 0B1;
    Q_filtered_10b[1097] = 086;
    Q_filtered_10b[1096] = 055;
    Q_filtered_10b[1095] = 01F;
    Q_filtered_10b[1094] = 3E4;
    Q_filtered_10b[1093] = 3AB;
    Q_filtered_10b[1092] = 37B;
    Q_filtered_10b[1091] = 34D;
    Q_filtered_10b[1090] = 32C;
    Q_filtered_10b[1089] = 317;
    Q_filtered_10b[1088] = 312;
    Q_filtered_10b[1087] = 315;
    Q_filtered_10b[1086] = 32A;
    Q_filtered_10b[1085] = 34B;
    Q_filtered_10b[1084] = 378;
    Q_filtered_10b[1083] = 3A9;
    Q_filtered_10b[1082] = 3E4;
    Q_filtered_10b[1081] = 023;
    Q_filtered_10b[1080] = 05C;
    Q_filtered_10b[1079] = 090;
    Q_filtered_10b[1078] = 0BA;
    Q_filtered_10b[1077] = 0DB;
    Q_filtered_10b[1076] = 0ED;
    Q_filtered_10b[1075] = 0EE;
    Q_filtered_10b[1074] = 0E4;
    Q_filtered_10b[1073] = 0CC;
    Q_filtered_10b[1072] = 0AB;
    Q_filtered_10b[1071] = 07E;
    Q_filtered_10b[1070] = 050;
    Q_filtered_10b[1069] = 01B;
    Q_filtered_10b[1068] = 3E8;
    Q_filtered_10b[1067] = 3B9;
    Q_filtered_10b[1066] = 38E;
    Q_filtered_10b[1065] = 36A;
    Q_filtered_10b[1064] = 34F;
    Q_filtered_10b[1063] = 33A;
    Q_filtered_10b[1062] = 333;
    Q_filtered_10b[1061] = 32E;
    Q_filtered_10b[1060] = 331;
    Q_filtered_10b[1059] = 33A;
    Q_filtered_10b[1058] = 349;
    Q_filtered_10b[1057] = 353;
    Q_filtered_10b[1056] = 363;
    Q_filtered_10b[1055] = 374;
    Q_filtered_10b[1054] = 37F;
    Q_filtered_10b[1053] = 38B;
    Q_filtered_10b[1052] = 392;
    Q_filtered_10b[1051] = 399;
    Q_filtered_10b[1050] = 39A;
    Q_filtered_10b[1049] = 398;
    Q_filtered_10b[1048] = 394;
    Q_filtered_10b[1047] = 38F;
    Q_filtered_10b[1046] = 388;
    Q_filtered_10b[1045] = 37F;
    Q_filtered_10b[1044] = 377;
    Q_filtered_10b[1043] = 36A;
    Q_filtered_10b[1042] = 35E;
    Q_filtered_10b[1041] = 356;
    Q_filtered_10b[1040] = 34D;
    Q_filtered_10b[1039] = 347;
    Q_filtered_10b[1038] = 342;
    Q_filtered_10b[1037] = 342;
    Q_filtered_10b[1036] = 349;
    Q_filtered_10b[1035] = 351;
    Q_filtered_10b[1034] = 35D;
    Q_filtered_10b[1033] = 368;
    Q_filtered_10b[1032] = 379;
    Q_filtered_10b[1031] = 386;
    Q_filtered_10b[1030] = 398;
    Q_filtered_10b[1029] = 3A5;
    Q_filtered_10b[1028] = 3B1;
    Q_filtered_10b[1027] = 3C1;
    Q_filtered_10b[1026] = 3C9;
    Q_filtered_10b[1025] = 3D2;
    Q_filtered_10b[1024] = 3DB;
    Q_filtered_10b[1023] = 3E4;
    Q_filtered_10b[1022] = 3EB;
    Q_filtered_10b[1021] = 3F7;
    Q_filtered_10b[1020] = 004;
    Q_filtered_10b[1019] = 014;
    Q_filtered_10b[1018] = 02A;
    Q_filtered_10b[1017] = 043;
    Q_filtered_10b[1016] = 05E;
    Q_filtered_10b[1015] = 07B;
    Q_filtered_10b[1014] = 096;
    Q_filtered_10b[1013] = 0AF;
    Q_filtered_10b[1012] = 0C2;
    Q_filtered_10b[1011] = 0CE;
    Q_filtered_10b[1010] = 0D2;
    Q_filtered_10b[1009] = 0CE;
    Q_filtered_10b[1008] = 0BF;
    Q_filtered_10b[1007] = 0A9;
    Q_filtered_10b[1006] = 08E;
    Q_filtered_10b[1005] = 06C;
    Q_filtered_10b[1004] = 049;
    Q_filtered_10b[1003] = 025;
    Q_filtered_10b[1002] = 003;
    Q_filtered_10b[1001] = 3E6;
    Q_filtered_10b[1000] = 3CE;
    Q_filtered_10b[999] = 3BC;
    Q_filtered_10b[998] = 3AD;
    Q_filtered_10b[997] = 3A5;
    Q_filtered_10b[996] = 39F;
    Q_filtered_10b[995] = 39C;
    Q_filtered_10b[994] = 39C;
    Q_filtered_10b[993] = 39E;
    Q_filtered_10b[992] = 39B;
    Q_filtered_10b[991] = 39A;
    Q_filtered_10b[990] = 398;
    Q_filtered_10b[989] = 394;
    Q_filtered_10b[988] = 38F;
    Q_filtered_10b[987] = 38B;
    Q_filtered_10b[986] = 388;
    Q_filtered_10b[985] = 384;
    Q_filtered_10b[984] = 382;
    Q_filtered_10b[983] = 383;
    Q_filtered_10b[982] = 385;
    Q_filtered_10b[981] = 389;
    Q_filtered_10b[980] = 38C;
    Q_filtered_10b[979] = 392;
    Q_filtered_10b[978] = 397;
    Q_filtered_10b[977] = 39B;
    Q_filtered_10b[976] = 39F;
    Q_filtered_10b[975] = 3A3;
    Q_filtered_10b[974] = 3A2;
    Q_filtered_10b[973] = 3A3;
    Q_filtered_10b[972] = 3A6;
    Q_filtered_10b[971] = 3AB;
    Q_filtered_10b[970] = 3B0;
    Q_filtered_10b[969] = 3BC;
    Q_filtered_10b[968] = 3CA;
    Q_filtered_10b[967] = 3DC;
    Q_filtered_10b[966] = 3F4;
    Q_filtered_10b[965] = 00D;
    Q_filtered_10b[964] = 028;
    Q_filtered_10b[963] = 045;
    Q_filtered_10b[962] = 05F;
    Q_filtered_10b[961] = 078;
    Q_filtered_10b[960] = 08B;
    Q_filtered_10b[959] = 099;
    Q_filtered_10b[958] = 09F;
    Q_filtered_10b[957] = 09F;
    Q_filtered_10b[956] = 095;
    Q_filtered_10b[955] = 082;
    Q_filtered_10b[954] = 06B;
    Q_filtered_10b[953] = 04D;
    Q_filtered_10b[952] = 02B;
    Q_filtered_10b[951] = 006;
    Q_filtered_10b[950] = 3E5;
    Q_filtered_10b[949] = 3C7;
    Q_filtered_10b[948] = 3B1;
    Q_filtered_10b[947] = 39F;
    Q_filtered_10b[946] = 395;
    Q_filtered_10b[945] = 395;
    Q_filtered_10b[944] = 39B;
    Q_filtered_10b[943] = 3A6;
    Q_filtered_10b[942] = 3B5;
    Q_filtered_10b[941] = 3CA;
    Q_filtered_10b[940] = 3DE;
    Q_filtered_10b[939] = 3F5;
    Q_filtered_10b[938] = 009;
    Q_filtered_10b[937] = 01A;
    Q_filtered_10b[936] = 02B;
    Q_filtered_10b[935] = 037;
    Q_filtered_10b[934] = 040;
    Q_filtered_10b[933] = 048;
    Q_filtered_10b[932] = 04A;
    Q_filtered_10b[931] = 04F;
    Q_filtered_10b[930] = 054;
    Q_filtered_10b[929] = 05A;
    Q_filtered_10b[928] = 05F;
    Q_filtered_10b[927] = 06B;
    Q_filtered_10b[926] = 077;
    Q_filtered_10b[925] = 085;
    Q_filtered_10b[924] = 094;
    Q_filtered_10b[923] = 0A1;
    Q_filtered_10b[922] = 0AD;
    Q_filtered_10b[921] = 0B6;
    Q_filtered_10b[920] = 0BC;
    Q_filtered_10b[919] = 0BC;
    Q_filtered_10b[918] = 0BA;
    Q_filtered_10b[917] = 0B1;
    Q_filtered_10b[916] = 0A5;
    Q_filtered_10b[915] = 095;
    Q_filtered_10b[914] = 083;
    Q_filtered_10b[913] = 071;
    Q_filtered_10b[912] = 05F;
    Q_filtered_10b[911] = 04D;
    Q_filtered_10b[910] = 03D;
    Q_filtered_10b[909] = 02F;
    Q_filtered_10b[908] = 025;
    Q_filtered_10b[907] = 01A;
    Q_filtered_10b[906] = 011;
    Q_filtered_10b[905] = 00A;
    Q_filtered_10b[904] = 002;
    Q_filtered_10b[903] = 3FD;
    Q_filtered_10b[902] = 3F7;
    Q_filtered_10b[901] = 3F0;
    Q_filtered_10b[900] = 3E6;
    Q_filtered_10b[899] = 3DF;
    Q_filtered_10b[898] = 3D7;
    Q_filtered_10b[897] = 3CC;
    Q_filtered_10b[896] = 3C6;
    Q_filtered_10b[895] = 3C0;
    Q_filtered_10b[894] = 3BA;
    Q_filtered_10b[893] = 3B6;
    Q_filtered_10b[892] = 3B4;
    Q_filtered_10b[891] = 3B1;
    Q_filtered_10b[890] = 3AE;
    Q_filtered_10b[889] = 3AA;
    Q_filtered_10b[888] = 3A4;
    Q_filtered_10b[887] = 39E;
    Q_filtered_10b[886] = 395;
    Q_filtered_10b[885] = 389;
    Q_filtered_10b[884] = 381;
    Q_filtered_10b[883] = 373;
    Q_filtered_10b[882] = 36A;
    Q_filtered_10b[881] = 366;
    Q_filtered_10b[880] = 367;
    Q_filtered_10b[879] = 36B;
    Q_filtered_10b[878] = 37C;
    Q_filtered_10b[877] = 393;
    Q_filtered_10b[876] = 3B1;
    Q_filtered_10b[875] = 3D8;
    Q_filtered_10b[874] = 004;
    Q_filtered_10b[873] = 035;
    Q_filtered_10b[872] = 064;
    Q_filtered_10b[871] = 08E;
    Q_filtered_10b[870] = 0B2;
    Q_filtered_10b[869] = 0CE;
    Q_filtered_10b[868] = 0DF;
    Q_filtered_10b[867] = 0E3;
    Q_filtered_10b[866] = 0DC;
    Q_filtered_10b[865] = 0C9;
    Q_filtered_10b[864] = 0AD;
    Q_filtered_10b[863] = 088;
    Q_filtered_10b[862] = 060;
    Q_filtered_10b[861] = 031;
    Q_filtered_10b[860] = 004;
    Q_filtered_10b[859] = 3DC;
    Q_filtered_10b[858] = 3B7;
    Q_filtered_10b[857] = 39C;
    Q_filtered_10b[856] = 387;
    Q_filtered_10b[855] = 377;
    Q_filtered_10b[854] = 372;
    Q_filtered_10b[853] = 36F;
    Q_filtered_10b[852] = 36E;
    Q_filtered_10b[851] = 36E;
    Q_filtered_10b[850] = 372;
    Q_filtered_10b[849] = 36D;
    Q_filtered_10b[848] = 36A;
    Q_filtered_10b[847] = 363;
    Q_filtered_10b[846] = 358;
    Q_filtered_10b[845] = 350;
    Q_filtered_10b[844] = 347;
    Q_filtered_10b[843] = 340;
    Q_filtered_10b[842] = 33D;
    Q_filtered_10b[841] = 33E;
    Q_filtered_10b[840] = 345;
    Q_filtered_10b[839] = 354;
    Q_filtered_10b[838] = 367;
    Q_filtered_10b[837] = 37E;
    Q_filtered_10b[836] = 39C;
    Q_filtered_10b[835] = 3BA;
    Q_filtered_10b[834] = 3D7;
    Q_filtered_10b[833] = 3F6;
    Q_filtered_10b[832] = 011;
    Q_filtered_10b[831] = 027;
    Q_filtered_10b[830] = 038;
    Q_filtered_10b[829] = 04A;
    Q_filtered_10b[828] = 055;
    Q_filtered_10b[827] = 05F;
    Q_filtered_10b[826] = 068;
    Q_filtered_10b[825] = 06C;
    Q_filtered_10b[824] = 070;
    Q_filtered_10b[823] = 077;
    Q_filtered_10b[822] = 07F;
    Q_filtered_10b[821] = 085;
    Q_filtered_10b[820] = 08E;
    Q_filtered_10b[819] = 098;
    Q_filtered_10b[818] = 0A1;
    Q_filtered_10b[817] = 0A8;
    Q_filtered_10b[816] = 0AE;
    Q_filtered_10b[815] = 0B1;
    Q_filtered_10b[814] = 0B2;
    Q_filtered_10b[813] = 0AF;
    Q_filtered_10b[812] = 0AB;
    Q_filtered_10b[811] = 0A7;
    Q_filtered_10b[810] = 0A1;
    Q_filtered_10b[809] = 09E;
    Q_filtered_10b[808] = 09C;
    Q_filtered_10b[807] = 099;
    Q_filtered_10b[806] = 098;
    Q_filtered_10b[805] = 097;
    Q_filtered_10b[804] = 097;
    Q_filtered_10b[803] = 091;
    Q_filtered_10b[802] = 089;
    Q_filtered_10b[801] = 07E;
    Q_filtered_10b[800] = 06C;
    Q_filtered_10b[799] = 05B;
    Q_filtered_10b[798] = 044;
    Q_filtered_10b[797] = 029;
    Q_filtered_10b[796] = 00D;
    Q_filtered_10b[795] = 3F4;
    Q_filtered_10b[794] = 3D8;
    Q_filtered_10b[793] = 3BE;
    Q_filtered_10b[792] = 3A6;
    Q_filtered_10b[791] = 395;
    Q_filtered_10b[790] = 383;
    Q_filtered_10b[789] = 377;
    Q_filtered_10b[788] = 36E;
    Q_filtered_10b[787] = 368;
    Q_filtered_10b[786] = 367;
    Q_filtered_10b[785] = 367;
    Q_filtered_10b[784] = 366;
    Q_filtered_10b[783] = 366;
    Q_filtered_10b[782] = 369;
    Q_filtered_10b[781] = 367;
    Q_filtered_10b[780] = 366;
    Q_filtered_10b[779] = 360;
    Q_filtered_10b[778] = 35D;
    Q_filtered_10b[777] = 357;
    Q_filtered_10b[776] = 354;
    Q_filtered_10b[775] = 350;
    Q_filtered_10b[774] = 350;
    Q_filtered_10b[773] = 353;
    Q_filtered_10b[772] = 357;
    Q_filtered_10b[771] = 35D;
    Q_filtered_10b[770] = 364;
    Q_filtered_10b[769] = 36D;
    Q_filtered_10b[768] = 376;
    Q_filtered_10b[767] = 37E;
    Q_filtered_10b[766] = 384;
    Q_filtered_10b[765] = 38A;
    Q_filtered_10b[764] = 38E;
    Q_filtered_10b[763] = 393;
    Q_filtered_10b[762] = 393;
    Q_filtered_10b[761] = 394;
    Q_filtered_10b[760] = 391;
    Q_filtered_10b[759] = 390;
    Q_filtered_10b[758] = 38B;
    Q_filtered_10b[757] = 386;
    Q_filtered_10b[756] = 37F;
    Q_filtered_10b[755] = 37C;
    Q_filtered_10b[754] = 379;
    Q_filtered_10b[753] = 379;
    Q_filtered_10b[752] = 378;
    Q_filtered_10b[751] = 37B;
    Q_filtered_10b[750] = 382;
    Q_filtered_10b[749] = 388;
    Q_filtered_10b[748] = 391;
    Q_filtered_10b[747] = 398;
    Q_filtered_10b[746] = 3A2;
    Q_filtered_10b[745] = 3AA;
    Q_filtered_10b[744] = 3B5;
    Q_filtered_10b[743] = 3BB;
    Q_filtered_10b[742] = 3C2;
    Q_filtered_10b[741] = 3CC;
    Q_filtered_10b[740] = 3D1;
    Q_filtered_10b[739] = 3D7;
    Q_filtered_10b[738] = 3DD;
    Q_filtered_10b[737] = 3E4;
    Q_filtered_10b[736] = 3E9;
    Q_filtered_10b[735] = 3F2;
    Q_filtered_10b[734] = 3FC;
    Q_filtered_10b[733] = 009;
    Q_filtered_10b[732] = 019;
    Q_filtered_10b[731] = 02B;
    Q_filtered_10b[730] = 03E;
    Q_filtered_10b[729] = 054;
    Q_filtered_10b[728] = 067;
    Q_filtered_10b[727] = 07B;
    Q_filtered_10b[726] = 08A;
    Q_filtered_10b[725] = 095;
    Q_filtered_10b[724] = 099;
    Q_filtered_10b[723] = 099;
    Q_filtered_10b[722] = 08F;
    Q_filtered_10b[721] = 07D;
    Q_filtered_10b[720] = 067;
    Q_filtered_10b[719] = 04B;
    Q_filtered_10b[718] = 02A;
    Q_filtered_10b[717] = 006;
    Q_filtered_10b[716] = 3E6;
    Q_filtered_10b[715] = 3C8;
    Q_filtered_10b[714] = 3B2;
    Q_filtered_10b[713] = 3A0;
    Q_filtered_10b[712] = 396;
    Q_filtered_10b[711] = 395;
    Q_filtered_10b[710] = 39A;
    Q_filtered_10b[709] = 3A5;
    Q_filtered_10b[708] = 3B4;
    Q_filtered_10b[707] = 3C9;
    Q_filtered_10b[706] = 3DD;
    Q_filtered_10b[705] = 3F5;
    Q_filtered_10b[704] = 00A;
    Q_filtered_10b[703] = 01B;
    Q_filtered_10b[702] = 02D;
    Q_filtered_10b[701] = 038;
    Q_filtered_10b[700] = 041;
    Q_filtered_10b[699] = 048;
    Q_filtered_10b[698] = 04A;
    Q_filtered_10b[697] = 04E;
    Q_filtered_10b[696] = 052;
    Q_filtered_10b[695] = 058;
    Q_filtered_10b[694] = 05D;
    Q_filtered_10b[693] = 06A;
    Q_filtered_10b[692] = 074;
    Q_filtered_10b[691] = 082;
    Q_filtered_10b[690] = 093;
    Q_filtered_10b[689] = 09E;
    Q_filtered_10b[688] = 0AE;
    Q_filtered_10b[687] = 0B8;
    Q_filtered_10b[686] = 0C0;
    Q_filtered_10b[685] = 0C2;
    Q_filtered_10b[684] = 0C2;
    Q_filtered_10b[683] = 0B8;
    Q_filtered_10b[682] = 0A8;
    Q_filtered_10b[681] = 093;
    Q_filtered_10b[680] = 079;
    Q_filtered_10b[679] = 05A;
    Q_filtered_10b[678] = 038;
    Q_filtered_10b[677] = 018;
    Q_filtered_10b[676] = 3FB;
    Q_filtered_10b[675] = 3E4;
    Q_filtered_10b[674] = 3D2;
    Q_filtered_10b[673] = 3C7;
    Q_filtered_10b[672] = 3C3;
    Q_filtered_10b[671] = 3C8;
    Q_filtered_10b[670] = 3D2;
    Q_filtered_10b[669] = 3E1;
    Q_filtered_10b[668] = 3F5;
    Q_filtered_10b[667] = 00B;
    Q_filtered_10b[666] = 023;
    Q_filtered_10b[665] = 03A;
    Q_filtered_10b[664] = 04D;
    Q_filtered_10b[663] = 05E;
    Q_filtered_10b[662] = 06B;
    Q_filtered_10b[661] = 075;
    Q_filtered_10b[660] = 07D;
    Q_filtered_10b[659] = 07E;
    Q_filtered_10b[658] = 082;
    Q_filtered_10b[657] = 084;
    Q_filtered_10b[656] = 086;
    Q_filtered_10b[655] = 086;
    Q_filtered_10b[654] = 08D;
    Q_filtered_10b[653] = 093;
    Q_filtered_10b[652] = 09A;
    Q_filtered_10b[651] = 0A2;
    Q_filtered_10b[650] = 0A8;
    Q_filtered_10b[649] = 0AD;
    Q_filtered_10b[648] = 0B1;
    Q_filtered_10b[647] = 0B3;
    Q_filtered_10b[646] = 0B1;
    Q_filtered_10b[645] = 0AE;
    Q_filtered_10b[644] = 0A7;
    Q_filtered_10b[643] = 0A0;
    Q_filtered_10b[642] = 097;
    Q_filtered_10b[641] = 08D;
    Q_filtered_10b[640] = 084;
    Q_filtered_10b[639] = 07D;
    Q_filtered_10b[638] = 075;
    Q_filtered_10b[637] = 06D;
    Q_filtered_10b[636] = 067;
    Q_filtered_10b[635] = 062;
    Q_filtered_10b[634] = 059;
    Q_filtered_10b[633] = 050;
    Q_filtered_10b[632] = 046;
    Q_filtered_10b[631] = 037;
    Q_filtered_10b[630] = 02A;
    Q_filtered_10b[629] = 019;
    Q_filtered_10b[628] = 005;
    Q_filtered_10b[627] = 3EF;
    Q_filtered_10b[626] = 3DC;
    Q_filtered_10b[625] = 3C6;
    Q_filtered_10b[624] = 3B1;
    Q_filtered_10b[623] = 39D;
    Q_filtered_10b[622] = 38F;
    Q_filtered_10b[621] = 380;
    Q_filtered_10b[620] = 377;
    Q_filtered_10b[619] = 371;
    Q_filtered_10b[618] = 36E;
    Q_filtered_10b[617] = 371;
    Q_filtered_10b[616] = 374;
    Q_filtered_10b[615] = 378;
    Q_filtered_10b[614] = 37C;
    Q_filtered_10b[613] = 382;
    Q_filtered_10b[612] = 385;
    Q_filtered_10b[611] = 387;
    Q_filtered_10b[610] = 387;
    Q_filtered_10b[609] = 388;
    Q_filtered_10b[608] = 387;
    Q_filtered_10b[607] = 388;
    Q_filtered_10b[606] = 388;
    Q_filtered_10b[605] = 38A;
    Q_filtered_10b[604] = 38D;
    Q_filtered_10b[603] = 390;
    Q_filtered_10b[602] = 394;
    Q_filtered_10b[601] = 398;
    Q_filtered_10b[600] = 39B;
    Q_filtered_10b[599] = 3A0;
    Q_filtered_10b[598] = 3A4;
    Q_filtered_10b[597] = 3A7;
    Q_filtered_10b[596] = 3AA;
    Q_filtered_10b[595] = 3AF;
    Q_filtered_10b[594] = 3B6;
    Q_filtered_10b[593] = 3BB;
    Q_filtered_10b[592] = 3C3;
    Q_filtered_10b[591] = 3C9;
    Q_filtered_10b[590] = 3D2;
    Q_filtered_10b[589] = 3DB;
    Q_filtered_10b[588] = 3E7;
    Q_filtered_10b[587] = 3F0;
    Q_filtered_10b[586] = 3FA;
    Q_filtered_10b[585] = 006;
    Q_filtered_10b[584] = 00C;
    Q_filtered_10b[583] = 013;
    Q_filtered_10b[582] = 018;
    Q_filtered_10b[581] = 01C;
    Q_filtered_10b[580] = 01D;
    Q_filtered_10b[579] = 01F;
    Q_filtered_10b[578] = 022;
    Q_filtered_10b[577] = 025;
    Q_filtered_10b[576] = 02B;
    Q_filtered_10b[575] = 032;
    Q_filtered_10b[574] = 03D;
    Q_filtered_10b[573] = 048;
    Q_filtered_10b[572] = 052;
    Q_filtered_10b[571] = 05D;
    Q_filtered_10b[570] = 065;
    Q_filtered_10b[569] = 067;
    Q_filtered_10b[568] = 066;
    Q_filtered_10b[567] = 05E;
    Q_filtered_10b[566] = 04E;
    Q_filtered_10b[565] = 03A;
    Q_filtered_10b[564] = 021;
    Q_filtered_10b[563] = 002;
    Q_filtered_10b[562] = 3E1;
    Q_filtered_10b[561] = 3C0;
    Q_filtered_10b[560] = 39E;
    Q_filtered_10b[559] = 381;
    Q_filtered_10b[558] = 368;
    Q_filtered_10b[557] = 355;
    Q_filtered_10b[556] = 345;
    Q_filtered_10b[555] = 33E;
    Q_filtered_10b[554] = 33A;
    Q_filtered_10b[553] = 33C;
    Q_filtered_10b[552] = 343;
    Q_filtered_10b[551] = 34D;
    Q_filtered_10b[550] = 356;
    Q_filtered_10b[549] = 362;
    Q_filtered_10b[548] = 36F;
    Q_filtered_10b[547] = 378;
    Q_filtered_10b[546] = 381;
    Q_filtered_10b[545] = 385;
    Q_filtered_10b[544] = 38A;
    Q_filtered_10b[543] = 38C;
    Q_filtered_10b[542] = 38D;
    Q_filtered_10b[541] = 38D;
    Q_filtered_10b[540] = 38F;
    Q_filtered_10b[539] = 390;
    Q_filtered_10b[538] = 392;
    Q_filtered_10b[537] = 396;
    Q_filtered_10b[536] = 39A;
    Q_filtered_10b[535] = 39F;
    Q_filtered_10b[534] = 3A5;
    Q_filtered_10b[533] = 3AC;
    Q_filtered_10b[532] = 3AF;
    Q_filtered_10b[531] = 3B3;
    Q_filtered_10b[530] = 3B6;
    Q_filtered_10b[529] = 3BB;
    Q_filtered_10b[528] = 3BC;
    Q_filtered_10b[527] = 3BF;
    Q_filtered_10b[526] = 3C1;
    Q_filtered_10b[525] = 3C6;
    Q_filtered_10b[524] = 3C9;
    Q_filtered_10b[523] = 3D0;
    Q_filtered_10b[522] = 3D8;
    Q_filtered_10b[521] = 3DF;
    Q_filtered_10b[520] = 3E9;
    Q_filtered_10b[519] = 3EF;
    Q_filtered_10b[518] = 3F6;
    Q_filtered_10b[517] = 3F8;
    Q_filtered_10b[516] = 3FA;
    Q_filtered_10b[515] = 3F5;
    Q_filtered_10b[514] = 3EE;
    Q_filtered_10b[513] = 3E5;
    Q_filtered_10b[512] = 3DA;
    Q_filtered_10b[511] = 3CC;
    Q_filtered_10b[510] = 3BC;
    Q_filtered_10b[509] = 3AD;
    Q_filtered_10b[508] = 3A1;
    Q_filtered_10b[507] = 395;
    Q_filtered_10b[506] = 390;
    Q_filtered_10b[505] = 38A;
    Q_filtered_10b[504] = 387;
    Q_filtered_10b[503] = 388;
    Q_filtered_10b[502] = 388;
    Q_filtered_10b[501] = 388;
    Q_filtered_10b[500] = 384;
    Q_filtered_10b[499] = 382;
    Q_filtered_10b[498] = 378;
    Q_filtered_10b[497] = 36F;
    Q_filtered_10b[496] = 360;
    Q_filtered_10b[495] = 351;
    Q_filtered_10b[494] = 346;
    Q_filtered_10b[493] = 339;
    Q_filtered_10b[492] = 330;
    Q_filtered_10b[491] = 32E;
    Q_filtered_10b[490] = 333;
    Q_filtered_10b[489] = 33D;
    Q_filtered_10b[488] = 353;
    Q_filtered_10b[487] = 36E;
    Q_filtered_10b[486] = 391;
    Q_filtered_10b[485] = 3BB;
    Q_filtered_10b[484] = 3EA;
    Q_filtered_10b[483] = 018;
    Q_filtered_10b[482] = 047;
    Q_filtered_10b[481] = 072;
    Q_filtered_10b[480] = 096;
    Q_filtered_10b[479] = 0B2;
    Q_filtered_10b[478] = 0C8;
    Q_filtered_10b[477] = 0D2;
    Q_filtered_10b[476] = 0D5;
    Q_filtered_10b[475] = 0D0;
    Q_filtered_10b[474] = 0C3;
    Q_filtered_10b[473] = 0B2;
    Q_filtered_10b[472] = 0A0;
    Q_filtered_10b[471] = 08C;
    Q_filtered_10b[470] = 077;
    Q_filtered_10b[469] = 068;
    Q_filtered_10b[468] = 05A;
    Q_filtered_10b[467] = 052;
    Q_filtered_10b[466] = 04B;
    Q_filtered_10b[465] = 046;
    Q_filtered_10b[464] = 045;
    Q_filtered_10b[463] = 043;
    Q_filtered_10b[462] = 03E;
    Q_filtered_10b[461] = 039;
    Q_filtered_10b[460] = 035;
    Q_filtered_10b[459] = 02A;
    Q_filtered_10b[458] = 020;
    Q_filtered_10b[457] = 014;
    Q_filtered_10b[456] = 007;
    Q_filtered_10b[455] = 3FB;
    Q_filtered_10b[454] = 3F2;
    Q_filtered_10b[453] = 3EB;
    Q_filtered_10b[452] = 3E4;
    Q_filtered_10b[451] = 3DE;
    Q_filtered_10b[450] = 3DD;
    Q_filtered_10b[449] = 3DC;
    Q_filtered_10b[448] = 3DD;
    Q_filtered_10b[447] = 3DE;
    Q_filtered_10b[446] = 3E1;
    Q_filtered_10b[445] = 3E2;
    Q_filtered_10b[444] = 3E4;
    Q_filtered_10b[443] = 3E4;
    Q_filtered_10b[442] = 3E3;
    Q_filtered_10b[441] = 3E0;
    Q_filtered_10b[440] = 3DF;
    Q_filtered_10b[439] = 3DE;
    Q_filtered_10b[438] = 3DE;
    Q_filtered_10b[437] = 3E1;
    Q_filtered_10b[436] = 3E6;
    Q_filtered_10b[435] = 3EE;
    Q_filtered_10b[434] = 3F7;
    Q_filtered_10b[433] = 004;
    Q_filtered_10b[432] = 010;
    Q_filtered_10b[431] = 01E;
    Q_filtered_10b[430] = 02C;
    Q_filtered_10b[429] = 038;
    Q_filtered_10b[428] = 043;
    Q_filtered_10b[427] = 04B;
    Q_filtered_10b[426] = 052;
    Q_filtered_10b[425] = 055;
    Q_filtered_10b[424] = 057;
    Q_filtered_10b[423] = 055;
    Q_filtered_10b[422] = 050;
    Q_filtered_10b[421] = 049;
    Q_filtered_10b[420] = 041;
    Q_filtered_10b[419] = 039;
    Q_filtered_10b[418] = 02F;
    Q_filtered_10b[417] = 025;
    Q_filtered_10b[416] = 01E;
    Q_filtered_10b[415] = 016;
    Q_filtered_10b[414] = 011;
    Q_filtered_10b[413] = 00D;
    Q_filtered_10b[412] = 00C;
    Q_filtered_10b[411] = 00C;
    Q_filtered_10b[410] = 00E;
    Q_filtered_10b[409] = 014;
    Q_filtered_10b[408] = 01B;
    Q_filtered_10b[407] = 023;
    Q_filtered_10b[406] = 02D;
    Q_filtered_10b[405] = 038;
    Q_filtered_10b[404] = 043;
    Q_filtered_10b[403] = 04B;
    Q_filtered_10b[402] = 054;
    Q_filtered_10b[401] = 05A;
    Q_filtered_10b[400] = 05D;
    Q_filtered_10b[399] = 05B;
    Q_filtered_10b[398] = 057;
    Q_filtered_10b[397] = 04E;
    Q_filtered_10b[396] = 042;
    Q_filtered_10b[395] = 031;
    Q_filtered_10b[394] = 01F;
    Q_filtered_10b[393] = 00A;
    Q_filtered_10b[392] = 3F5;
    Q_filtered_10b[391] = 3E0;
    Q_filtered_10b[390] = 3CD;
    Q_filtered_10b[389] = 3BB;
    Q_filtered_10b[388] = 3AE;
    Q_filtered_10b[387] = 3A4;
    Q_filtered_10b[386] = 3A0;
    Q_filtered_10b[385] = 39F;
    Q_filtered_10b[384] = 3A4;
    Q_filtered_10b[383] = 3AE;
    Q_filtered_10b[382] = 3BB;
    Q_filtered_10b[381] = 3CB;
    Q_filtered_10b[380] = 3DB;
    Q_filtered_10b[379] = 3ED;
    Q_filtered_10b[378] = 3FE;
    Q_filtered_10b[377] = 00C;
    Q_filtered_10b[376] = 01A;
    Q_filtered_10b[375] = 024;
    Q_filtered_10b[374] = 02B;
    Q_filtered_10b[373] = 02D;
    Q_filtered_10b[372] = 02E;
    Q_filtered_10b[371] = 029;
    Q_filtered_10b[370] = 01F;
    Q_filtered_10b[369] = 012;
    Q_filtered_10b[368] = 002;
    Q_filtered_10b[367] = 3EF;
    Q_filtered_10b[366] = 3D8;
    Q_filtered_10b[365] = 3C4;
    Q_filtered_10b[364] = 3B1;
    Q_filtered_10b[363] = 3A2;
    Q_filtered_10b[362] = 396;
    Q_filtered_10b[361] = 392;
    Q_filtered_10b[360] = 395;
    Q_filtered_10b[359] = 39E;
    Q_filtered_10b[358] = 3AF;
    Q_filtered_10b[357] = 3C4;
    Q_filtered_10b[356] = 3E0;
    Q_filtered_10b[355] = 3FF;
    Q_filtered_10b[354] = 023;
    Q_filtered_10b[353] = 045;
    Q_filtered_10b[352] = 066;
    Q_filtered_10b[351] = 085;
    Q_filtered_10b[350] = 09D;
    Q_filtered_10b[349] = 0B0;
    Q_filtered_10b[348] = 0BE;
    Q_filtered_10b[347] = 0C2;
    Q_filtered_10b[346] = 0C3;
    Q_filtered_10b[345] = 0BF;
    Q_filtered_10b[344] = 0B8;
    Q_filtered_10b[343] = 0AD;
    Q_filtered_10b[342] = 0A6;
    Q_filtered_10b[341] = 09D;
    Q_filtered_10b[340] = 098;
    Q_filtered_10b[339] = 094;
    Q_filtered_10b[338] = 090;
    Q_filtered_10b[337] = 08E;
    Q_filtered_10b[336] = 08C;
    Q_filtered_10b[335] = 088;
    Q_filtered_10b[334] = 083;
    Q_filtered_10b[333] = 07B;
    Q_filtered_10b[332] = 06E;
    Q_filtered_10b[331] = 061;
    Q_filtered_10b[330] = 050;
    Q_filtered_10b[329] = 03B;
    Q_filtered_10b[328] = 026;
    Q_filtered_10b[327] = 013;
    Q_filtered_10b[326] = 3FC;
    Q_filtered_10b[325] = 3E9;
    Q_filtered_10b[324] = 3D7;
    Q_filtered_10b[323] = 3CA;
    Q_filtered_10b[322] = 3BB;
    Q_filtered_10b[321] = 3B0;
    Q_filtered_10b[320] = 3A6;
    Q_filtered_10b[319] = 39D;
    Q_filtered_10b[318] = 398;
    Q_filtered_10b[317] = 392;
    Q_filtered_10b[316] = 38A;
    Q_filtered_10b[315] = 383;
    Q_filtered_10b[314] = 37F;
    Q_filtered_10b[313] = 376;
    Q_filtered_10b[312] = 36E;
    Q_filtered_10b[311] = 363;
    Q_filtered_10b[310] = 35C;
    Q_filtered_10b[309] = 353;
    Q_filtered_10b[308] = 34F;
    Q_filtered_10b[307] = 34A;
    Q_filtered_10b[306] = 34A;
    Q_filtered_10b[305] = 34E;
    Q_filtered_10b[304] = 353;
    Q_filtered_10b[303] = 35B;
    Q_filtered_10b[302] = 362;
    Q_filtered_10b[301] = 36C;
    Q_filtered_10b[300] = 376;
    Q_filtered_10b[299] = 37E;
    Q_filtered_10b[298] = 385;
    Q_filtered_10b[297] = 38A;
    Q_filtered_10b[296] = 38E;
    Q_filtered_10b[295] = 393;
    Q_filtered_10b[294] = 393;
    Q_filtered_10b[293] = 394;
    Q_filtered_10b[292] = 392;
    Q_filtered_10b[291] = 390;
    Q_filtered_10b[290] = 38B;
    Q_filtered_10b[289] = 385;
    Q_filtered_10b[288] = 37D;
    Q_filtered_10b[287] = 378;
    Q_filtered_10b[286] = 374;
    Q_filtered_10b[285] = 373;
    Q_filtered_10b[284] = 371;
    Q_filtered_10b[283] = 375;
    Q_filtered_10b[282] = 37D;
    Q_filtered_10b[281] = 385;
    Q_filtered_10b[280] = 392;
    Q_filtered_10b[279] = 39C;
    Q_filtered_10b[278] = 3AC;
    Q_filtered_10b[277] = 3B9;
    Q_filtered_10b[276] = 3CB;
    Q_filtered_10b[275] = 3D8;
    Q_filtered_10b[274] = 3E5;
    Q_filtered_10b[273] = 3F5;
    Q_filtered_10b[272] = 3FE;
    Q_filtered_10b[271] = 007;
    Q_filtered_10b[270] = 010;
    Q_filtered_10b[269] = 017;
    Q_filtered_10b[268] = 01C;
    Q_filtered_10b[267] = 025;
    Q_filtered_10b[266] = 02E;
    Q_filtered_10b[265] = 03A;
    Q_filtered_10b[264] = 04B;
    Q_filtered_10b[263] = 05E;
    Q_filtered_10b[262] = 074;
    Q_filtered_10b[261] = 08C;
    Q_filtered_10b[260] = 0A2;
    Q_filtered_10b[259] = 0B7;
    Q_filtered_10b[258] = 0C7;
    Q_filtered_10b[257] = 0D1;
    Q_filtered_10b[256] = 0D2;
    Q_filtered_10b[255] = 0CC;
    Q_filtered_10b[254] = 0BB;
    Q_filtered_10b[253] = 0A2;
    Q_filtered_10b[252] = 082;
    Q_filtered_10b[251] = 05B;
    Q_filtered_10b[250] = 032;
    Q_filtered_10b[249] = 008;
    Q_filtered_10b[248] = 3DE;
    Q_filtered_10b[247] = 3BA;
    Q_filtered_10b[246] = 39B;
    Q_filtered_10b[245] = 383;
    Q_filtered_10b[244] = 370;
    Q_filtered_10b[243] = 367;
    Q_filtered_10b[242] = 361;
    Q_filtered_10b[241] = 363;
    Q_filtered_10b[240] = 36B;
    Q_filtered_10b[239] = 378;
    Q_filtered_10b[238] = 383;
    Q_filtered_10b[237] = 392;
    Q_filtered_10b[236] = 3A3;
    Q_filtered_10b[235] = 3AF;
    Q_filtered_10b[234] = 3BA;
    Q_filtered_10b[233] = 3C1;
    Q_filtered_10b[232] = 3C7;
    Q_filtered_10b[231] = 3C8;
    Q_filtered_10b[230] = 3C6;
    Q_filtered_10b[229] = 3C2;
    Q_filtered_10b[228] = 3BD;
    Q_filtered_10b[227] = 3B7;
    Q_filtered_10b[226] = 3AE;
    Q_filtered_10b[225] = 3A7;
    Q_filtered_10b[224] = 39E;
    Q_filtered_10b[223] = 395;
    Q_filtered_10b[222] = 38E;
    Q_filtered_10b[221] = 387;
    Q_filtered_10b[220] = 380;
    Q_filtered_10b[219] = 37C;
    Q_filtered_10b[218] = 37A;
    Q_filtered_10b[217] = 37D;
    Q_filtered_10b[216] = 37F;
    Q_filtered_10b[215] = 386;
    Q_filtered_10b[214] = 38D;
    Q_filtered_10b[213] = 399;
    Q_filtered_10b[212] = 3A3;
    Q_filtered_10b[211] = 3B1;
    Q_filtered_10b[210] = 3BD;
    Q_filtered_10b[209] = 3CA;
    Q_filtered_10b[208] = 3D7;
    Q_filtered_10b[207] = 3E1;
    Q_filtered_10b[206] = 3E9;
    Q_filtered_10b[205] = 3F0;
    Q_filtered_10b[204] = 3F4;
    Q_filtered_10b[203] = 3F5;
    Q_filtered_10b[202] = 3F6;
    Q_filtered_10b[201] = 3F3;
    Q_filtered_10b[200] = 3F1;
    Q_filtered_10b[199] = 3EE;
    Q_filtered_10b[198] = 3EB;
    Q_filtered_10b[197] = 3E8;
    Q_filtered_10b[196] = 3E7;
    Q_filtered_10b[195] = 3E7;
    Q_filtered_10b[194] = 3E6;
    Q_filtered_10b[193] = 3E7;
    Q_filtered_10b[192] = 3E7;
    Q_filtered_10b[191] = 3E9;
    Q_filtered_10b[190] = 3E9;
    Q_filtered_10b[189] = 3E9;
    Q_filtered_10b[188] = 3E9;
    Q_filtered_10b[187] = 3EA;
    Q_filtered_10b[186] = 3E9;
    Q_filtered_10b[185] = 3EA;
    Q_filtered_10b[184] = 3EB;
    Q_filtered_10b[183] = 3EB;
    Q_filtered_10b[182] = 3ED;
    Q_filtered_10b[181] = 3EE;
    Q_filtered_10b[180] = 3F0;
    Q_filtered_10b[179] = 3EF;
    Q_filtered_10b[178] = 3EF;
    Q_filtered_10b[177] = 3EC;
    Q_filtered_10b[176] = 3E8;
    Q_filtered_10b[175] = 3E4;
    Q_filtered_10b[174] = 3DF;
    Q_filtered_10b[173] = 3D8;
    Q_filtered_10b[172] = 3D3;
    Q_filtered_10b[171] = 3CE;
    Q_filtered_10b[170] = 3C8;
    Q_filtered_10b[169] = 3C4;
    Q_filtered_10b[168] = 3BE;
    Q_filtered_10b[167] = 3BB;
    Q_filtered_10b[166] = 3B7;
    Q_filtered_10b[165] = 3B6;
    Q_filtered_10b[164] = 3B2;
    Q_filtered_10b[163] = 3B1;
    Q_filtered_10b[162] = 3B1;
    Q_filtered_10b[161] = 3B2;
    Q_filtered_10b[160] = 3B3;
    Q_filtered_10b[159] = 3B5;
    Q_filtered_10b[158] = 3B9;
    Q_filtered_10b[157] = 3BC;
    Q_filtered_10b[156] = 3BF;
    Q_filtered_10b[155] = 3C0;
    Q_filtered_10b[154] = 3C2;
    Q_filtered_10b[153] = 3C1;
    Q_filtered_10b[152] = 3C1;
    Q_filtered_10b[151] = 3BC;
    Q_filtered_10b[150] = 3B8;
    Q_filtered_10b[149] = 3B3;
    Q_filtered_10b[148] = 3AE;
    Q_filtered_10b[147] = 3A7;
    Q_filtered_10b[146] = 39F;
    Q_filtered_10b[145] = 398;
    Q_filtered_10b[144] = 392;
    Q_filtered_10b[143] = 38D;
    Q_filtered_10b[142] = 38A;
    Q_filtered_10b[141] = 387;
    Q_filtered_10b[140] = 386;
    Q_filtered_10b[139] = 388;
    Q_filtered_10b[138] = 388;
    Q_filtered_10b[137] = 38A;
    Q_filtered_10b[136] = 389;
    Q_filtered_10b[135] = 38A;
    Q_filtered_10b[134] = 387;
    Q_filtered_10b[133] = 385;
    Q_filtered_10b[132] = 37F;
    Q_filtered_10b[131] = 37A;
    Q_filtered_10b[130] = 377;
    Q_filtered_10b[129] = 373;
    Q_filtered_10b[128] = 370;
    Q_filtered_10b[127] = 372;
    Q_filtered_10b[126] = 377;
    Q_filtered_10b[125] = 37E;
    Q_filtered_10b[124] = 38C;
    Q_filtered_10b[123] = 39A;
    Q_filtered_10b[122] = 3AE;
    Q_filtered_10b[121] = 3C4;
    Q_filtered_10b[120] = 3DE;
    Q_filtered_10b[119] = 3F6;
    Q_filtered_10b[118] = 00F;
    Q_filtered_10b[117] = 027;
    Q_filtered_10b[116] = 039;
    Q_filtered_10b[115] = 048;
    Q_filtered_10b[114] = 054;
    Q_filtered_10b[113] = 05B;
    Q_filtered_10b[112] = 05C;
    Q_filtered_10b[111] = 05C;
    Q_filtered_10b[110] = 059;
    Q_filtered_10b[109] = 055;
    Q_filtered_10b[108] = 053;
    Q_filtered_10b[107] = 050;
    Q_filtered_10b[106] = 04F;
    Q_filtered_10b[105] = 051;
    Q_filtered_10b[104] = 052;
    Q_filtered_10b[103] = 057;
    Q_filtered_10b[102] = 05A;
    Q_filtered_10b[101] = 05B;
    Q_filtered_10b[100] = 05B;
    Q_filtered_10b[99] = 056;
    Q_filtered_10b[98] = 04B;
    Q_filtered_10b[97] = 03C;
    Q_filtered_10b[96] = 02A;
    Q_filtered_10b[95] = 011;
    Q_filtered_10b[94] = 3F5;
    Q_filtered_10b[93] = 3D8;
    Q_filtered_10b[92] = 3BB;
    Q_filtered_10b[91] = 3A1;
    Q_filtered_10b[90] = 38C;
    Q_filtered_10b[89] = 37C;
    Q_filtered_10b[88] = 370;
    Q_filtered_10b[87] = 36C;
    Q_filtered_10b[86] = 36E;
    Q_filtered_10b[85] = 374;
    Q_filtered_10b[84] = 37F;
    Q_filtered_10b[83] = 38D;
    Q_filtered_10b[82] = 39B;
    Q_filtered_10b[81] = 3AA;
    Q_filtered_10b[80] = 3B7;
    Q_filtered_10b[79] = 3C2;
    Q_filtered_10b[78] = 3CC;
    Q_filtered_10b[77] = 3D3;
    Q_filtered_10b[76] = 3D9;
    Q_filtered_10b[75] = 3DF;
    Q_filtered_10b[74] = 3E4;
    Q_filtered_10b[73] = 3EB;
    Q_filtered_10b[72] = 3F4;
    Q_filtered_10b[71] = 3FE;
    Q_filtered_10b[70] = 009;
    Q_filtered_10b[69] = 019;
    Q_filtered_10b[68] = 02A;
    Q_filtered_10b[67] = 03A;
    Q_filtered_10b[66] = 04C;
    Q_filtered_10b[65] = 05C;
    Q_filtered_10b[64] = 069;
    Q_filtered_10b[63] = 074;
    Q_filtered_10b[62] = 07E;
    Q_filtered_10b[61] = 083;
    Q_filtered_10b[60] = 087;
    Q_filtered_10b[59] = 088;
    Q_filtered_10b[58] = 086;
    Q_filtered_10b[57] = 084;
    Q_filtered_10b[56] = 083;
    Q_filtered_10b[55] = 081;
    Q_filtered_10b[54] = 080;
    Q_filtered_10b[53] = 080;
    Q_filtered_10b[52] = 080;
    Q_filtered_10b[51] = 084;
    Q_filtered_10b[50] = 085;
    Q_filtered_10b[49] = 086;
    Q_filtered_10b[48] = 083;
    Q_filtered_10b[47] = 080;
    Q_filtered_10b[46] = 078;
    Q_filtered_10b[45] = 06D;
    Q_filtered_10b[44] = 05F;
    Q_filtered_10b[43] = 04E;
    Q_filtered_10b[42] = 03C;
    Q_filtered_10b[41] = 029;
    Q_filtered_10b[40] = 014;
    Q_filtered_10b[39] = 002;
    Q_filtered_10b[38] = 3F3;
    Q_filtered_10b[37] = 3E7;
    Q_filtered_10b[36] = 3DC;
    Q_filtered_10b[35] = 3D6;
    Q_filtered_10b[34] = 3D4;
    Q_filtered_10b[33] = 3D4;
    Q_filtered_10b[32] = 3D9;
    Q_filtered_10b[31] = 3DE;
    Q_filtered_10b[30] = 3E5;
    Q_filtered_10b[29] = 3ED;
    Q_filtered_10b[28] = 3F5;
    Q_filtered_10b[27] = 3FB;
    Q_filtered_10b[26] = 000;
    Q_filtered_10b[25] = 002;
    Q_filtered_10b[24] = 004;
    Q_filtered_10b[23] = 004;
    Q_filtered_10b[22] = 003;
    Q_filtered_10b[21] = 002;
    Q_filtered_10b[20] = 000;
    Q_filtered_10b[19] = 000;
    Q_filtered_10b[18] = 3FE;
    Q_filtered_10b[17] = 3FF;
    Q_filtered_10b[16] = 3FE;
    Q_filtered_10b[15] = 3FF;
    Q_filtered_10b[14] = 000;
    Q_filtered_10b[13] = 3FF;
    Q_filtered_10b[12] = 3FF;
    Q_filtered_10b[11] = 3FF;
    Q_filtered_10b[10] = 000;
    Q_filtered_10b[9] = 000;
    Q_filtered_10b[8] = 000;
    Q_filtered_10b[7] = 000;
    Q_filtered_10b[6] = 000;
    Q_filtered_10b[5] = 001;
    Q_filtered_10b[4] = 000;
    Q_filtered_10b[3] = 000;
    Q_filtered_10b[2] = 000;
    Q_filtered_10b[1] = 000;
    Q_filtered_10b[0] = 000;


// I Channel 12b Expected output
//     first 64 samples only
    I_filtered_12b[63] = 000;
    I_filtered_12b[62] = 000;
    I_filtered_12b[61] = 005;
    I_filtered_12b[60] = 00A;
    I_filtered_12b[59] = 00A;
    I_filtered_12b[58] = 00F;
    I_filtered_12b[57] = 00A;
    I_filtered_12b[56] = 00A;
    I_filtered_12b[55] = 005;
    I_filtered_12b[54] = 000;
    I_filtered_12b[53] = FF6;
    I_filtered_12b[52] = FF1;
    I_filtered_12b[51] = FF1;
    I_filtered_12b[50] = FF1;
    I_filtered_12b[49] = FF6;
    I_filtered_12b[48] = FFA;
    I_filtered_12b[47] = 008;
    I_filtered_12b[46] = 017;
    I_filtered_12b[45] = 025;
    I_filtered_12b[44] = 035;
    I_filtered_12b[43] = 03F;
    I_filtered_12b[42] = 040;
    I_filtered_12b[41] = 03C;
    I_filtered_12b[40] = 02F;
    I_filtered_12b[39] = 00D;
    I_filtered_12b[38] = FE0;
    I_filtered_12b[37] = FA9;
    I_filtered_12b[36] = F62;
    I_filtered_12b[35] = F10;
    I_filtered_12b[34] = EBC;
    I_filtered_12b[33] = E64;
    I_filtered_12b[32] = E15;
    I_filtered_12b[31] = DD2;
    I_filtered_12b[30] = D9E;
    I_filtered_12b[29] = D81;
    I_filtered_12b[28] = D79;
    I_filtered_12b[27] = D88;
    I_filtered_12b[26] = DAE;
    I_filtered_12b[25] = DE9;
    I_filtered_12b[24] = E35;
    I_filtered_12b[23] = E8D;
    I_filtered_12b[22] = EEE;
    I_filtered_12b[21] = F48;
    I_filtered_12b[20] = FA6;
    I_filtered_12b[19] = FF5;
    I_filtered_12b[18] = 039;
    I_filtered_12b[17] = 06E;
    I_filtered_12b[16] = 09A;
    I_filtered_12b[15] = 0AF;
    I_filtered_12b[14] = 0BB;
    I_filtered_12b[13] = 0BF;
    I_filtered_12b[12] = 0B4;
    I_filtered_12b[11] = 0A3;
    I_filtered_12b[10] = 090;
    I_filtered_12b[9] = 082;
    I_filtered_12b[8] = 06F;
    I_filtered_12b[7] = 062;
    I_filtered_12b[6] = 05A;
    I_filtered_12b[5] = 04E;
    I_filtered_12b[4] = 049;
    I_filtered_12b[3] = 048;
    I_filtered_12b[2] = 04F;
    I_filtered_12b[1] = 050;
    I_filtered_12b[0] = 05F;


// Q Channel 12b Expected output
//     first 64 samples only
    Q_filtered_12b[63] = 000;
    Q_filtered_12b[62] = 000;
    Q_filtered_12b[61] = 001;
    Q_filtered_12b[60] = 002;
    Q_filtered_12b[59] = 002;
    Q_filtered_12b[58] = 003;
    Q_filtered_12b[57] = 002;
    Q_filtered_12b[56] = 002;
    Q_filtered_12b[55] = 001;
    Q_filtered_12b[54] = 000;
    Q_filtered_12b[53] = FFE;
    Q_filtered_12b[52] = FFD;
    Q_filtered_12b[51] = FFD;
    Q_filtered_12b[50] = FFD;
    Q_filtered_12b[49] = FFE;
    Q_filtered_12b[48] = FFA;
    Q_filtered_12b[47] = FF8;
    Q_filtered_12b[46] = FFB;
    Q_filtered_12b[45] = FF8;
    Q_filtered_12b[44] = 000;
    Q_filtered_12b[43] = 002;
    Q_filtered_12b[42] = 007;
    Q_filtered_12b[41] = 00B;
    Q_filtered_12b[40] = 012;
    Q_filtered_12b[39] = 011;
    Q_filtered_12b[38] = 009;
    Q_filtered_12b[37] = FFF;
    Q_filtered_12b[36] = FED;
    Q_filtered_12b[35] = FD5;
    Q_filtered_12b[34] = FB2;
    Q_filtered_12b[33] = F94;
    Q_filtered_12b[32] = F78;
    Q_filtered_12b[31] = F62;
    Q_filtered_12b[30] = F4F;
    Q_filtered_12b[29] = F4E;
    Q_filtered_12b[28] = F57;
    Q_filtered_12b[27] = F71;
    Q_filtered_12b[26] = F9A;
    Q_filtered_12b[25] = FCB;
    Q_filtered_12b[24] = 009;
    Q_filtered_12b[23] = 052;
    Q_filtered_12b[22] = 0A3;
    Q_filtered_12b[21] = 0EF;
    Q_filtered_12b[20] = 139;
    Q_filtered_12b[19] = 17E;
    Q_filtered_12b[18] = 1B4;
    Q_filtered_12b[17] = 1DF;
    Q_filtered_12b[16] = 202;
    Q_filtered_12b[15] = 20E;
    Q_filtered_12b[14] = 217;
    Q_filtered_12b[13] = 216;
    Q_filtered_12b[12] = 20F;
    Q_filtered_12b[11] = 202;
    Q_filtered_12b[10] = 201;
    Q_filtered_12b[9] = 1FF;
    Q_filtered_12b[8] = 204;
    Q_filtered_12b[7] = 20B;
    Q_filtered_12b[6] = 211;
    Q_filtered_12b[5] = 219;
    Q_filtered_12b[4] = 220;
    Q_filtered_12b[3] = 21C;
    Q_filtered_12b[2] = 20E;
    Q_filtered_12b[1] = 1F8;
    Q_filtered_12b[0] = 1D0;
end

endmodule

