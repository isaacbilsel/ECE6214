`timescale 1ns / 1ps
`include "modulator_signals.vh"

module baseband_dsp_tb;

    reg data_in;
    reg data_clk;
    reg dsp_clk;
    reg rst_n_data;
    reg rst_n_dsp;
    reg msg_in;
    reg rw;
    reg [9:0] mem_addr;
    reg [7:0] coeff_in; 
    reg enable;
    reg [3:0] sample_rate;
    reg mapping;
    wire mem_read_out;
    wire [9:0] I_out;
    wire [9:0] Q_out;

    baseband_dsp DUT(
        .data_in(data_in),
        .data_clk(data_clk),
        .dsp_clk(dsp_clk),
        .rst_n_data(rst_n_data),
        .rst_n_dsp(rst_n_dsp),
        .msg_in(msg_in),
        .rw(rw),
        .mem_addr(mem_addr),
        .coeff_in(coeff_in),
        .mem_read_out(mem_read_out),
        .I_out(I_out),
	    .Q_out(Q_out)
    );
	
	// Datastream variables
	reg [7:0] Icoeff [0:70];
	reg [7:0] Qcoeff [0:70];
	reg [779:0] datastream;
	reg [9:0] I_filtered_10b[0:1733];
	reg [9:0] Q_filtered_10b[0:1733];
	reg [11:0] I_filtered_12b[0:63]; //11
	reg [11:0] Q_filtered_12b[0:63]; //11
	
    always #8.333 data_clk = ~data_clk;
    always #3.846 dsp_clk = ~dsp_clk;
    
    reg [8*39:0] testcase;
    integer i;
	
    initial begin
        testcase = "Initializing";
        data_clk <= 1'b0;
        dsp_clk <= 1'b0;
        rst_n_data <= 1'b0;
        rst_n_dsp <= 1'b0;
		sample_rate <= 4'd13;
        data_in <= 1'b0; 
        enable <= 1'b0;

		repeat(2) @(posedge data_clk);
		rst_n_data <= 1'b1;
        enable <= 1'b1;
		@(posedge data_clk);

        @(posedge dsp_clk)
        rst_n_dsp <= 1'b1;
        @(posedge dsp_clk)

        // Write I coefficients to memory
        @(negedge dsp_clk);
		for (i=0; i<=70; i=i+1) begin
			msg_in <= 1'b1;
			rw <= 1'b1;
			mem_addr  <= i + 128;
			coeff_in  <= Icoeff[i];
			@(negedge dsp_clk);	 
		end

		// Write Q coefficients to memory
		for (i=0; i<=70; i = i+1) begin
			msg_in <= 1'b1;
			rw <= 1'b1;
			mem_addr  <= i + 256;
			coeff_in  <= Qcoeff[i];
			@(negedge dsp_clk);	 
		end
		msg_in <= 1'b0;

        testcase = "Coeff_Read";
        repeat(3) @(posedge dsp_clk);
        // Test reading coeff I memory
		// coeff_read_out should set to 0xFD
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr  <= 133; // This is addr of 5th I coeff: oxFD
		repeat(2) @(posedge dsp_clk);
		msg_in <= 1'b0;

		repeat(3) @(posedge dsp_clk);
		// Test reading coeff Q memory
		// coeff_read_out should set to 0x02
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr  <= 266; 
		repeat(3) @(posedge dsp_clk);
		msg_in <= 1'b0;

		// flush the pipeline
		repeat(5) @(posedge dsp_clk);

        // Send in datastream with 12 bit header
        testcase <= "Datastream";    
        @(negedge data_clk);
        for (i=779; i>=0; i=i-1) begin
            data_in <= datastream[i]; 
            @(negedge data_clk);
        end

        repeat(3) @(posedge dsp_clk);
        // Test reading I output memory
		// Should read 10th output: 0x00 or 0x05F idk
        testcase <= "Output_read"; 
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr <= 512;
		// Read last 4 LSBs
		repeat(1) @(posedge dsp_clk);
		mem_addr  <= 513;
		repeat(3) @(posedge dsp_clk);

		// Test reading I output memory
		// Should read 10th output: 0x090 or 0x082 or 0xFF6 idk
        testcase <= "Output_read"; 
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr <= 532;
		// Read last 4 LSBs
		repeat(1) @(posedge dsp_clk);
		mem_addr  <= 533;
		repeat(3) @(posedge dsp_clk);

        // Write compare outputs function and log file
        $finish;
    end

initial begin
    // I filter coefficients
    Icoeff[0] = 8'h00;
    Icoeff[1] = 8'h00;
    Icoeff[2] = 8'hFF;
    Icoeff[3] = 8'hFE;
    Icoeff[4] = 8'hFE;
    Icoeff[5] = 8'hFD;
    Icoeff[6] = 8'hFE;
    Icoeff[7] = 8'hFE;
    Icoeff[8] = 8'hFF;
    Icoeff[9] = 8'h00;
    Icoeff[10] = 8'h02;
    Icoeff[11] = 8'h03;
    Icoeff[12] = 8'h03;
    Icoeff[13] = 8'h03;
    Icoeff[14] = 8'h02;
    Icoeff[15] = 8'h01;
    Icoeff[16] = 8'hFE;
    Icoeff[17] = 8'hFB;
    Icoeff[18] = 8'hF8;
    Icoeff[19] = 8'hF5;
    Icoeff[20] = 8'hF3;
    Icoeff[21] = 8'hF3;
    Icoeff[22] = 8'hF4;
    Icoeff[23] = 8'hF7;
    Icoeff[24] = 8'hFE;
    Icoeff[25] = 8'h07;
    Icoeff[26] = 8'h12;
    Icoeff[27] = 8'h20;
    Icoeff[28] = 8'h30;
    Icoeff[29] = 8'h40;
    Icoeff[30] = 8'h51;
    Icoeff[31] = 8'h60;
    Icoeff[32] = 8'h6D;
    Icoeff[33] = 8'h77;
    Icoeff[34] = 8'h7D;
    Icoeff[35] = 8'h7F;
    Icoeff[36] = 8'h7D;
    Icoeff[37] = 8'h77;
    Icoeff[38] = 8'h6D;
    Icoeff[39] = 8'h60;
    Icoeff[40] = 8'h51;
    Icoeff[41] = 8'h40;
    Icoeff[42] = 8'h30;
    Icoeff[43] = 8'h20;
    Icoeff[44] = 8'h12;
    Icoeff[45] = 8'h07;
    Icoeff[46] = 8'hFE;
    Icoeff[47] = 8'hF7;
    Icoeff[48] = 8'hF4;
    Icoeff[49] = 8'hF3;
    Icoeff[50] = 8'hF3;
    Icoeff[51] = 8'hF5;
    Icoeff[52] = 8'hF8;
    Icoeff[53] = 8'hFB;
    Icoeff[54] = 8'hFE;
    Icoeff[55] = 8'h01;
    Icoeff[56] = 8'h02;
    Icoeff[57] = 8'h03;
    Icoeff[58] = 8'h03;
    Icoeff[59] = 8'h03;
    Icoeff[60] = 8'h02;
    Icoeff[61] = 8'h00;
    Icoeff[62] = 8'hFF;
    Icoeff[63] = 8'hFE;
    Icoeff[64] = 8'hFE;
    Icoeff[65] = 8'hFD;
    Icoeff[66] = 8'hFE;
    Icoeff[67] = 8'hFE;
    Icoeff[68] = 8'hFF;
    Icoeff[69] = 8'h00;
    Icoeff[70] = 8'h00;


// Q filter coefficients
    Qcoeff[0] = 8'h00;
    Qcoeff[1] = 8'h00;
    Qcoeff[2] = 8'hFF;
    Qcoeff[3] = 8'hFE;
    Qcoeff[4] = 8'hFE;
    Qcoeff[5] = 8'hFD;
    Qcoeff[6] = 8'hFE;
    Qcoeff[7] = 8'hFE;
    Qcoeff[8] = 8'hFF;
    Qcoeff[9] = 8'h00;
    Qcoeff[10] = 8'h02;
    Qcoeff[11] = 8'h03;
    Qcoeff[12] = 8'h03;
    Qcoeff[13] = 8'h03;
    Qcoeff[14] = 8'h02;
    Qcoeff[15] = 8'h01;
    Qcoeff[16] = 8'hFE;
    Qcoeff[17] = 8'hFB;
    Qcoeff[18] = 8'hF9;
    Qcoeff[19] = 8'hF6;
    Qcoeff[20] = 8'hF4;
    Qcoeff[21] = 8'hF4;
    Qcoeff[22] = 8'hF5;
    Qcoeff[23] = 8'hF8;
    Qcoeff[24] = 8'hFE;
    Qcoeff[25] = 8'h06;
    Qcoeff[26] = 8'h10;
    Qcoeff[27] = 8'h1D;
    Qcoeff[28] = 8'h2B;
    Qcoeff[29] = 8'h3A;
    Qcoeff[30] = 8'h49;
    Qcoeff[31] = 8'h56;
    Qcoeff[32] = 8'h62;
    Qcoeff[33] = 8'h6B;
    Qcoeff[34] = 8'h71;
    Qcoeff[35] = 8'h72;
    Qcoeff[36] = 8'h71;
    Qcoeff[37] = 8'h6B;
    Qcoeff[38] = 8'h62;
    Qcoeff[39] = 8'h56;
    Qcoeff[40] = 8'h49;
    Qcoeff[41] = 8'h3A;
    Qcoeff[42] = 8'h2B;
    Qcoeff[43] = 8'h1D;
    Qcoeff[44] = 8'h10;
    Qcoeff[45] = 8'h06;
    Qcoeff[46] = 8'hFE;
    Qcoeff[47] = 8'hF8;
    Qcoeff[48] = 8'hF5;
    Qcoeff[49] = 8'hF4;
    Qcoeff[50] = 8'hF4;
    Qcoeff[51] = 8'hF6;
    Qcoeff[52] = 8'hF9;
    Qcoeff[53] = 8'hFB;
    Qcoeff[54] = 8'hFE;
    Qcoeff[55] = 8'h01;
    Qcoeff[56] = 8'h02;
    Qcoeff[57] = 8'h03;
    Qcoeff[58] = 8'h03;
    Qcoeff[59] = 8'h03;
    Qcoeff[60] = 8'h02;
    Qcoeff[61] = 8'h00;
    Qcoeff[62] = 8'hFF;
    Qcoeff[63] = 8'hFE;
    Qcoeff[64] = 8'hFE;
    Qcoeff[65] = 8'hFD;
    Qcoeff[66] = 8'hFE;
    Qcoeff[67] = 8'hFE;
    Qcoeff[68] = 8'hFF;
    Qcoeff[69] = 8'h00;
    Qcoeff[70] = 8'h00;


// Transmit Datastream with header
    [779:768] datastream = 12'hB38;
    [767:752] datastream = 16'hD196;
    [751:736] datastream = 16'h7592;
    [735:720] datastream = 16'hFAE7;
    [719:704] datastream = 16'h8104;
    [703:688] datastream = 16'h35D3;
    [687:672] datastream = 16'h6897;
    [671:656] datastream = 16'h9BF2;
    [655:640] datastream = 16'hA590;
    [639:624] datastream = 16'h451B;
    [623:608] datastream = 16'hE113;
    [607:592] datastream = 16'h15AC;
    [591:576] datastream = 16'hCB73;
    [575:560] datastream = 16'hDEBF;
    [559:544] datastream = 16'h0193;
    [543:528] datastream = 16'h6465;
    [527:512] datastream = 16'h02F3;
    [511:496] datastream = 16'h9786;
    [495:480] datastream = 16'h4A79;
    [479:464] datastream = 16'h6B6F;
    [463:448] datastream = 16'h2E55;
    [447:432] datastream = 16'hCDA6;
    [431:416] datastream = 16'h8028;
    [415:400] datastream = 16'h5FE6;
    [399:384] datastream = 16'h80E7;
    [383:368] datastream = 16'hFE45;
    [367:352] datastream = 16'h8CF6;
    [351:336] datastream = 16'hC49A;
    [335:320] datastream = 16'h4E25;
    [319:304] datastream = 16'hF8C8;
    [303:288] datastream = 16'h0985;
    [287:272] datastream = 16'hFC5F;
    [271:256] datastream = 16'h23B5;
    [255:240] datastream = 16'h94F7;
    [239:224] datastream = 16'hB931;
    [223:208] datastream = 16'hE1FA;
    [207:192] datastream = 16'h6604;
    [191:176] datastream = 16'hCB9A;
    [175:160] datastream = 16'hEA5C;
    [159:144] datastream = 16'h2DE4;
    [143:128] datastream = 16'hF7BA;
    [127:112] datastream = 16'h962F;
    [111:96] datastream = 16'h329D;
    [95:80] datastream = 16'h7727;
    [79:64] datastream = 16'h9533;
    [63:48] datastream = 16'h2149;
    [47:32] datastream = 16'h386A;
    [31:16] datastream = 16'hE179;
    [15:0] datastream = 16'hAA26;


// I Channel 10b Expected output
    I_filtered_10b[1733] = 10'h000;
    I_filtered_10b[1732] = 10'h000;
    I_filtered_10b[1731] = 10'h000;
    I_filtered_10b[1730] = 10'h000;
    I_filtered_10b[1729] = 10'h000;
    I_filtered_10b[1728] = 10'h000;
    I_filtered_10b[1727] = 10'h000;
    I_filtered_10b[1726] = 10'h000;
    I_filtered_10b[1725] = 10'h000;
    I_filtered_10b[1724] = 10'h000;
    I_filtered_10b[1723] = 10'h000;
    I_filtered_10b[1722] = 10'h000;
    I_filtered_10b[1721] = 10'h000;
    I_filtered_10b[1720] = 10'h000;
    I_filtered_10b[1719] = 10'h000;
    I_filtered_10b[1718] = 10'h000;
    I_filtered_10b[1717] = 10'h000;
    I_filtered_10b[1716] = 10'h001;
    I_filtered_10b[1715] = 10'h000;
    I_filtered_10b[1714] = 10'h000;
    I_filtered_10b[1713] = 10'h000;
    I_filtered_10b[1712] = 10'h000;
    I_filtered_10b[1711] = 10'h000;
    I_filtered_10b[1710] = 10'h3FF;
    I_filtered_10b[1709] = 10'h3FF;
    I_filtered_10b[1708] = 10'h3FF;
    I_filtered_10b[1707] = 10'h000;
    I_filtered_10b[1706] = 10'h001;
    I_filtered_10b[1705] = 10'h004;
    I_filtered_10b[1704] = 10'h005;
    I_filtered_10b[1703] = 10'h007;
    I_filtered_10b[1702] = 10'h006;
    I_filtered_10b[1701] = 10'h007;
    I_filtered_10b[1700] = 10'h005;
    I_filtered_10b[1699] = 10'h003;
    I_filtered_10b[1698] = 10'h3FF;
    I_filtered_10b[1697] = 10'h3FB;
    I_filtered_10b[1696] = 10'h3F9;
    I_filtered_10b[1695] = 10'h3F6;
    I_filtered_10b[1694] = 10'h3F5;
    I_filtered_10b[1693] = 10'h3F3;
    I_filtered_10b[1692] = 10'h3F5;
    I_filtered_10b[1691] = 10'h3F6;
    I_filtered_10b[1690] = 10'h3F8;
    I_filtered_10b[1689] = 10'h3FA;
    I_filtered_10b[1688] = 10'h3FB;
    I_filtered_10b[1687] = 10'h3F8;
    I_filtered_10b[1686] = 10'h3F5;
    I_filtered_10b[1685] = 10'h3EF;
    I_filtered_10b[1684] = 10'h3E4;
    I_filtered_10b[1683] = 10'h3D6;
    I_filtered_10b[1682] = 10'h3C6;
    I_filtered_10b[1681] = 10'h3B2;
    I_filtered_10b[1680] = 10'h39C;
    I_filtered_10b[1679] = 10'h386;
    I_filtered_10b[1678] = 10'h36F;
    I_filtered_10b[1677] = 10'h35A;
    I_filtered_10b[1676] = 10'h348;
    I_filtered_10b[1675] = 10'h33B;
    I_filtered_10b[1674] = 10'h332;
    I_filtered_10b[1673] = 10'h32E;
    I_filtered_10b[1672] = 10'h32F;
    I_filtered_10b[1671] = 10'h334;
    I_filtered_10b[1670] = 10'h33E;
    I_filtered_10b[1669] = 10'h34C;
    I_filtered_10b[1668] = 10'h35B;
    I_filtered_10b[1667] = 10'h36C;
    I_filtered_10b[1666] = 10'h37C;
    I_filtered_10b[1665] = 10'h38C;
    I_filtered_10b[1664] = 10'h399;
    I_filtered_10b[1663] = 10'h3A4;
    I_filtered_10b[1662] = 10'h3AC;
    I_filtered_10b[1661] = 10'h3B5;
    I_filtered_10b[1660] = 10'h3B9;
    I_filtered_10b[1659] = 10'h3BC;
    I_filtered_10b[1658] = 10'h3BF;
    I_filtered_10b[1657] = 10'h3C1;
    I_filtered_10b[1656] = 10'h3C3;
    I_filtered_10b[1655] = 10'h3C5;
    I_filtered_10b[1654] = 10'h3C7;
    I_filtered_10b[1653] = 10'h3C8;
    I_filtered_10b[1652] = 10'h3CD;
    I_filtered_10b[1651] = 10'h3D0;
    I_filtered_10b[1650] = 10'h3D5;
    I_filtered_10b[1649] = 10'h3D9;
    I_filtered_10b[1648] = 10'h3E0;
    I_filtered_10b[1647] = 10'h3E6;
    I_filtered_10b[1646] = 10'h3ED;
    I_filtered_10b[1645] = 10'h3F3;
    I_filtered_10b[1644] = 10'h3F6;
    I_filtered_10b[1643] = 10'h3FC;
    I_filtered_10b[1642] = 10'h3FE;
    I_filtered_10b[1641] = 10'h002;
    I_filtered_10b[1640] = 10'h003;
    I_filtered_10b[1639] = 10'h005;
    I_filtered_10b[1638] = 10'h008;
    I_filtered_10b[1637] = 10'h00A;
    I_filtered_10b[1636] = 10'h00C;
    I_filtered_10b[1635] = 10'h010;
    I_filtered_10b[1634] = 10'h014;
    I_filtered_10b[1633] = 10'h017;
    I_filtered_10b[1632] = 10'h01F;
    I_filtered_10b[1631] = 10'h027;
    I_filtered_10b[1630] = 10'h032;
    I_filtered_10b[1629] = 10'h03E;
    I_filtered_10b[1628] = 10'h04E;
    I_filtered_10b[1627] = 10'h05D;
    I_filtered_10b[1626] = 10'h06E;
    I_filtered_10b[1625] = 10'h07E;
    I_filtered_10b[1624] = 10'h08C;
    I_filtered_10b[1623] = 10'h097;
    I_filtered_10b[1622] = 10'h09D;
    I_filtered_10b[1621] = 10'h09F;
    I_filtered_10b[1620] = 10'h09B;
    I_filtered_10b[1619] = 10'h092;
    I_filtered_10b[1618] = 10'h083;
    I_filtered_10b[1617] = 10'h071;
    I_filtered_10b[1616] = 10'h05C;
    I_filtered_10b[1615] = 10'h043;
    I_filtered_10b[1614] = 10'h02C;
    I_filtered_10b[1613] = 10'h015;
    I_filtered_10b[1612] = 10'h000;
    I_filtered_10b[1611] = 10'h3F1;
    I_filtered_10b[1610] = 10'h3E3;
    I_filtered_10b[1609] = 10'h3D9;
    I_filtered_10b[1608] = 10'h3D4;
    I_filtered_10b[1607] = 10'h3D3;
    I_filtered_10b[1606] = 10'h3D3;
    I_filtered_10b[1605] = 10'h3D6;
    I_filtered_10b[1604] = 10'h3DA;
    I_filtered_10b[1603] = 10'h3DE;
    I_filtered_10b[1602] = 10'h3E1;
    I_filtered_10b[1601] = 10'h3E3;
    I_filtered_10b[1600] = 10'h3E4;
    I_filtered_10b[1599] = 10'h3E3;
    I_filtered_10b[1598] = 10'h3E3;
    I_filtered_10b[1597] = 10'h3E2;
    I_filtered_10b[1596] = 10'h3E2;
    I_filtered_10b[1595] = 10'h3E0;
    I_filtered_10b[1594] = 10'h3E2;
    I_filtered_10b[1593] = 10'h3E5;
    I_filtered_10b[1592] = 10'h3E9;
    I_filtered_10b[1591] = 10'h3ED;
    I_filtered_10b[1590] = 10'h3F4;
    I_filtered_10b[1589] = 10'h3FC;
    I_filtered_10b[1588] = 10'h002;
    I_filtered_10b[1587] = 10'h009;
    I_filtered_10b[1586] = 10'h00F;
    I_filtered_10b[1585] = 10'h012;
    I_filtered_10b[1584] = 10'h015;
    I_filtered_10b[1583] = 10'h018;
    I_filtered_10b[1582] = 10'h01A;
    I_filtered_10b[1581] = 10'h01A;
    I_filtered_10b[1580] = 10'h01E;
    I_filtered_10b[1579] = 10'h021;
    I_filtered_10b[1578] = 10'h026;
    I_filtered_10b[1577] = 10'h02C;
    I_filtered_10b[1576] = 10'h035;
    I_filtered_10b[1575] = 10'h040;
    I_filtered_10b[1574] = 10'h04A;
    I_filtered_10b[1573] = 10'h055;
    I_filtered_10b[1572] = 10'h05D;
    I_filtered_10b[1571] = 10'h064;
    I_filtered_10b[1570] = 10'h066;
    I_filtered_10b[1569] = 10'h065;
    I_filtered_10b[1568] = 10'h05F;
    I_filtered_10b[1567] = 10'h054;
    I_filtered_10b[1566] = 10'h046;
    I_filtered_10b[1565] = 10'h035;
    I_filtered_10b[1564] = 10'h021;
    I_filtered_10b[1563] = 10'h00A;
    I_filtered_10b[1562] = 10'h3F6;
    I_filtered_10b[1561] = 10'h3E1;
    I_filtered_10b[1560] = 10'h3CE;
    I_filtered_10b[1559] = 10'h3C1;
    I_filtered_10b[1558] = 10'h3B5;
    I_filtered_10b[1557] = 10'h3AC;
    I_filtered_10b[1556] = 10'h3A7;
    I_filtered_10b[1555] = 10'h3A5;
    I_filtered_10b[1554] = 10'h3A1;
    I_filtered_10b[1553] = 10'h39F;
    I_filtered_10b[1552] = 10'h39D;
    I_filtered_10b[1551] = 10'h399;
    I_filtered_10b[1550] = 10'h393;
    I_filtered_10b[1549] = 10'h38C;
    I_filtered_10b[1548] = 10'h381;
    I_filtered_10b[1547] = 10'h378;
    I_filtered_10b[1546] = 10'h36D;
    I_filtered_10b[1545] = 10'h366;
    I_filtered_10b[1544] = 10'h363;
    I_filtered_10b[1543] = 10'h361;
    I_filtered_10b[1542] = 10'h366;
    I_filtered_10b[1541] = 10'h371;
    I_filtered_10b[1540] = 10'h383;
    I_filtered_10b[1539] = 10'h399;
    I_filtered_10b[1538] = 10'h3B5;
    I_filtered_10b[1537] = 10'h3D5;
    I_filtered_10b[1536] = 10'h3F5;
    I_filtered_10b[1535] = 10'h016;
    I_filtered_10b[1534] = 10'h033;
    I_filtered_10b[1533] = 10'h04B;
    I_filtered_10b[1532] = 10'h05E;
    I_filtered_10b[1531] = 10'h06B;
    I_filtered_10b[1530] = 10'h071;
    I_filtered_10b[1529] = 10'h06F;
    I_filtered_10b[1528] = 10'h069;
    I_filtered_10b[1527] = 10'h05D;
    I_filtered_10b[1526] = 10'h04D;
    I_filtered_10b[1525] = 10'h03B;
    I_filtered_10b[1524] = 10'h026;
    I_filtered_10b[1523] = 10'h013;
    I_filtered_10b[1522] = 10'h003;
    I_filtered_10b[1521] = 10'h3F6;
    I_filtered_10b[1520] = 10'h3ED;
    I_filtered_10b[1519] = 10'h3E5;
    I_filtered_10b[1518] = 10'h3E1;
    I_filtered_10b[1517] = 10'h3E0;
    I_filtered_10b[1516] = 10'h3E1;
    I_filtered_10b[1515] = 10'h3DF;
    I_filtered_10b[1514] = 10'h3DC;
    I_filtered_10b[1513] = 10'h3DB;
    I_filtered_10b[1512] = 10'h3D4;
    I_filtered_10b[1511] = 10'h3CD;
    I_filtered_10b[1510] = 10'h3C3;
    I_filtered_10b[1509] = 10'h3B8;
    I_filtered_10b[1508] = 10'h3AE;
    I_filtered_10b[1507] = 10'h3A5;
    I_filtered_10b[1506] = 10'h39E;
    I_filtered_10b[1505] = 10'h39C;
    I_filtered_10b[1504] = 10'h39B;
    I_filtered_10b[1503] = 10'h3A0;
    I_filtered_10b[1502] = 10'h3A9;
    I_filtered_10b[1501] = 10'h3B7;
    I_filtered_10b[1500] = 10'h3C8;
    I_filtered_10b[1499] = 10'h3DD;
    I_filtered_10b[1498] = 10'h3F5;
    I_filtered_10b[1497] = 10'h00B;
    I_filtered_10b[1496] = 10'h022;
    I_filtered_10b[1495] = 10'h036;
    I_filtered_10b[1494] = 10'h045;
    I_filtered_10b[1493] = 10'h052;
    I_filtered_10b[1492] = 10'h05B;
    I_filtered_10b[1491] = 10'h05F;
    I_filtered_10b[1490] = 10'h05F;
    I_filtered_10b[1489] = 10'h060;
    I_filtered_10b[1488] = 10'h05D;
    I_filtered_10b[1487] = 10'h05A;
    I_filtered_10b[1486] = 10'h057;
    I_filtered_10b[1485] = 10'h054;
    I_filtered_10b[1484] = 10'h052;
    I_filtered_10b[1483] = 10'h054;
    I_filtered_10b[1482] = 10'h055;
    I_filtered_10b[1481] = 10'h05A;
    I_filtered_10b[1480] = 10'h05D;
    I_filtered_10b[1479] = 10'h05E;
    I_filtered_10b[1478] = 10'h05F;
    I_filtered_10b[1477] = 10'h05E;
    I_filtered_10b[1476] = 10'h056;
    I_filtered_10b[1475] = 10'h049;
    I_filtered_10b[1474] = 10'h03A;
    I_filtered_10b[1473] = 10'h025;
    I_filtered_10b[1472] = 10'h00C;
    I_filtered_10b[1471] = 10'h3F1;
    I_filtered_10b[1470] = 10'h3D4;
    I_filtered_10b[1469] = 10'h3BA;
    I_filtered_10b[1468] = 10'h3A6;
    I_filtered_10b[1467] = 10'h395;
    I_filtered_10b[1466] = 10'h38C;
    I_filtered_10b[1465] = 10'h389;
    I_filtered_10b[1464] = 10'h38F;
    I_filtered_10b[1463] = 10'h39D;
    I_filtered_10b[1462] = 10'h3B1;
    I_filtered_10b[1461] = 10'h3CA;
    I_filtered_10b[1460] = 10'h3E9;
    I_filtered_10b[1459] = 10'h00A;
    I_filtered_10b[1458] = 10'h02A;
    I_filtered_10b[1457] = 10'h049;
    I_filtered_10b[1456] = 10'h063;
    I_filtered_10b[1455] = 10'h078;
    I_filtered_10b[1454] = 10'h089;
    I_filtered_10b[1453] = 10'h094;
    I_filtered_10b[1452] = 10'h099;
    I_filtered_10b[1451] = 10'h099;
    I_filtered_10b[1450] = 10'h09A;
    I_filtered_10b[1449] = 10'h097;
    I_filtered_10b[1448] = 10'h091;
    I_filtered_10b[1447] = 10'h08F;
    I_filtered_10b[1446] = 10'h08C;
    I_filtered_10b[1445] = 10'h08C;
    I_filtered_10b[1444] = 10'h08E;
    I_filtered_10b[1443] = 10'h090;
    I_filtered_10b[1442] = 10'h093;
    I_filtered_10b[1441] = 10'h095;
    I_filtered_10b[1440] = 10'h093;
    I_filtered_10b[1439] = 10'h093;
    I_filtered_10b[1438] = 10'h08D;
    I_filtered_10b[1437] = 10'h084;
    I_filtered_10b[1436] = 10'h078;
    I_filtered_10b[1435] = 10'h069;
    I_filtered_10b[1434] = 10'h057;
    I_filtered_10b[1433] = 10'h041;
    I_filtered_10b[1432] = 10'h02D;
    I_filtered_10b[1431] = 10'h017;
    I_filtered_10b[1430] = 10'h004;
    I_filtered_10b[1429] = 10'h3F7;
    I_filtered_10b[1428] = 10'h3EB;
    I_filtered_10b[1427] = 10'h3E1;
    I_filtered_10b[1426] = 10'h3DA;
    I_filtered_10b[1425] = 10'h3D9;
    I_filtered_10b[1424] = 10'h3D5;
    I_filtered_10b[1423] = 10'h3D3;
    I_filtered_10b[1422] = 10'h3D1;
    I_filtered_10b[1421] = 10'h3CE;
    I_filtered_10b[1420] = 10'h3C8;
    I_filtered_10b[1419] = 10'h3C0;
    I_filtered_10b[1418] = 10'h3B6;
    I_filtered_10b[1417] = 10'h3AB;
    I_filtered_10b[1416] = 10'h3A1;
    I_filtered_10b[1415] = 10'h399;
    I_filtered_10b[1414] = 10'h396;
    I_filtered_10b[1413] = 10'h395;
    I_filtered_10b[1412] = 10'h39B;
    I_filtered_10b[1411] = 10'h3A7;
    I_filtered_10b[1410] = 10'h3BA;
    I_filtered_10b[1409] = 10'h3CF;
    I_filtered_10b[1408] = 10'h3EC;
    I_filtered_10b[1407] = 10'h00C;
    I_filtered_10b[1406] = 10'h02B;
    I_filtered_10b[1405] = 10'h04B;
    I_filtered_10b[1404] = 10'h067;
    I_filtered_10b[1403] = 10'h07C;
    I_filtered_10b[1402] = 10'h08E;
    I_filtered_10b[1401] = 10'h09A;
    I_filtered_10b[1400] = 10'h09F;
    I_filtered_10b[1399] = 10'h09D;
    I_filtered_10b[1398] = 10'h09A;
    I_filtered_10b[1397] = 10'h092;
    I_filtered_10b[1396] = 10'h088;
    I_filtered_10b[1395] = 10'h07F;
    I_filtered_10b[1394] = 10'h073;
    I_filtered_10b[1393] = 10'h06A;
    I_filtered_10b[1392] = 10'h066;
    I_filtered_10b[1391] = 10'h061;
    I_filtered_10b[1390] = 10'h062;
    I_filtered_10b[1389] = 10'h061;
    I_filtered_10b[1388] = 10'h05F;
    I_filtered_10b[1387] = 10'h05F;
    I_filtered_10b[1386] = 10'h05D;
    I_filtered_10b[1385] = 10'h052;
    I_filtered_10b[1384] = 10'h042;
    I_filtered_10b[1383] = 10'h02F;
    I_filtered_10b[1382] = 10'h013;
    I_filtered_10b[1381] = 10'h3F6;
    I_filtered_10b[1380] = 10'h3D4;
    I_filtered_10b[1379] = 10'h3AE;
    I_filtered_10b[1378] = 10'h38E;
    I_filtered_10b[1377] = 10'h36F;
    I_filtered_10b[1376] = 10'h358;
    I_filtered_10b[1375] = 10'h34A;
    I_filtered_10b[1374] = 10'h343;
    I_filtered_10b[1373] = 10'h348;
    I_filtered_10b[1372] = 10'h359;
    I_filtered_10b[1371] = 10'h377;
    I_filtered_10b[1370] = 10'h39C;
    I_filtered_10b[1369] = 10'h3CB;
    I_filtered_10b[1368] = 10'h3FE;
    I_filtered_10b[1367] = 10'h031;
    I_filtered_10b[1366] = 10'h067;
    I_filtered_10b[1365] = 10'h094;
    I_filtered_10b[1364] = 10'h0BD;
    I_filtered_10b[1363] = 10'h0DB;
    I_filtered_10b[1362] = 10'h0EF;
    I_filtered_10b[1361] = 10'h0F6;
    I_filtered_10b[1360] = 10'h0F4;
    I_filtered_10b[1359] = 10'h0E6;
    I_filtered_10b[1358] = 10'h0CB;
    I_filtered_10b[1357] = 10'h0A7;
    I_filtered_10b[1356] = 10'h07E;
    I_filtered_10b[1355] = 10'h04F;
    I_filtered_10b[1354] = 10'h020;
    I_filtered_10b[1353] = 10'h3F2;
    I_filtered_10b[1352] = 10'h3C8;
    I_filtered_10b[1351] = 10'h3A5;
    I_filtered_10b[1350] = 10'h38A;
    I_filtered_10b[1349] = 10'h37A;
    I_filtered_10b[1348] = 10'h377;
    I_filtered_10b[1347] = 10'h37C;
    I_filtered_10b[1346] = 10'h38D;
    I_filtered_10b[1345] = 10'h3A8;
    I_filtered_10b[1344] = 10'h3CB;
    I_filtered_10b[1343] = 10'h3F4;
    I_filtered_10b[1342] = 10'h021;
    I_filtered_10b[1341] = 10'h04E;
    I_filtered_10b[1340] = 10'h07A;
    I_filtered_10b[1339] = 10'h0A2;
    I_filtered_10b[1338] = 10'h0C4;
    I_filtered_10b[1337] = 10'h0DE;
    I_filtered_10b[1336] = 10'h0ED;
    I_filtered_10b[1335] = 10'h0F0;
    I_filtered_10b[1334] = 10'h0EC;
    I_filtered_10b[1333] = 10'h0DC;
    I_filtered_10b[1332] = 10'h0C2;
    I_filtered_10b[1331] = 10'h09F;
    I_filtered_10b[1330] = 10'h078;
    I_filtered_10b[1329] = 10'h04B;
    I_filtered_10b[1328] = 10'h01E;
    I_filtered_10b[1327] = 10'h3F3;
    I_filtered_10b[1326] = 10'h3CB;
    I_filtered_10b[1325] = 10'h3AA;
    I_filtered_10b[1324] = 10'h390;
    I_filtered_10b[1323] = 10'h381;
    I_filtered_10b[1322] = 10'h37D;
    I_filtered_10b[1321] = 10'h382;
    I_filtered_10b[1320] = 10'h390;
    I_filtered_10b[1319] = 10'h3A6;
    I_filtered_10b[1318] = 10'h3C4;
    I_filtered_10b[1317] = 10'h3E5;
    I_filtered_10b[1316] = 10'h00B;
    I_filtered_10b[1315] = 10'h02F;
    I_filtered_10b[1314] = 10'h051;
    I_filtered_10b[1313] = 10'h070;
    I_filtered_10b[1312] = 10'h087;
    I_filtered_10b[1311] = 10'h09A;
    I_filtered_10b[1310] = 10'h0A4;
    I_filtered_10b[1309] = 10'h0A5;
    I_filtered_10b[1308] = 10'h0A0;
    I_filtered_10b[1307] = 10'h098;
    I_filtered_10b[1306] = 10'h08C;
    I_filtered_10b[1305] = 10'h07B;
    I_filtered_10b[1304] = 10'h06C;
    I_filtered_10b[1303] = 10'h05A;
    I_filtered_10b[1302] = 10'h04D;
    I_filtered_10b[1301] = 10'h041;
    I_filtered_10b[1300] = 10'h036;
    I_filtered_10b[1299] = 10'h02C;
    I_filtered_10b[1298] = 10'h025;
    I_filtered_10b[1297] = 10'h01D;
    I_filtered_10b[1296] = 10'h01A;
    I_filtered_10b[1295] = 10'h014;
    I_filtered_10b[1294] = 10'h00D;
    I_filtered_10b[1293] = 10'h006;
    I_filtered_10b[1292] = 10'h3FF;
    I_filtered_10b[1291] = 10'h3F5;
    I_filtered_10b[1290] = 10'h3EC;
    I_filtered_10b[1289] = 10'h3E4;
    I_filtered_10b[1288] = 10'h3D8;
    I_filtered_10b[1287] = 10'h3D0;
    I_filtered_10b[1286] = 10'h3C5;
    I_filtered_10b[1285] = 10'h3BE;
    I_filtered_10b[1284] = 10'h3B5;
    I_filtered_10b[1283] = 10'h3AD;
    I_filtered_10b[1282] = 10'h3A6;
    I_filtered_10b[1281] = 10'h39E;
    I_filtered_10b[1280] = 10'h39B;
    I_filtered_10b[1279] = 10'h397;
    I_filtered_10b[1278] = 10'h394;
    I_filtered_10b[1277] = 10'h390;
    I_filtered_10b[1276] = 10'h38F;
    I_filtered_10b[1275] = 10'h38D;
    I_filtered_10b[1274] = 10'h38A;
    I_filtered_10b[1273] = 10'h387;
    I_filtered_10b[1272] = 10'h385;
    I_filtered_10b[1271] = 10'h382;
    I_filtered_10b[1270] = 10'h37F;
    I_filtered_10b[1269] = 10'h37D;
    I_filtered_10b[1268] = 10'h377;
    I_filtered_10b[1267] = 10'h373;
    I_filtered_10b[1266] = 10'h36D;
    I_filtered_10b[1265] = 10'h366;
    I_filtered_10b[1264] = 10'h35D;
    I_filtered_10b[1263] = 10'h354;
    I_filtered_10b[1262] = 10'h34B;
    I_filtered_10b[1261] = 10'h342;
    I_filtered_10b[1260] = 10'h33A;
    I_filtered_10b[1259] = 10'h334;
    I_filtered_10b[1258] = 10'h333;
    I_filtered_10b[1257] = 10'h334;
    I_filtered_10b[1256] = 10'h338;
    I_filtered_10b[1255] = 10'h341;
    I_filtered_10b[1254] = 10'h34E;
    I_filtered_10b[1253] = 10'h35F;
    I_filtered_10b[1252] = 10'h372;
    I_filtered_10b[1251] = 10'h388;
    I_filtered_10b[1250] = 10'h39C;
    I_filtered_10b[1249] = 10'h3B2;
    I_filtered_10b[1248] = 10'h3C6;
    I_filtered_10b[1247] = 10'h3D7;
    I_filtered_10b[1246] = 10'h3E5;
    I_filtered_10b[1245] = 10'h3F1;
    I_filtered_10b[1244] = 10'h3F8;
    I_filtered_10b[1243] = 10'h3FC;
    I_filtered_10b[1242] = 10'h3FD;
    I_filtered_10b[1241] = 10'h3FA;
    I_filtered_10b[1240] = 10'h3F6;
    I_filtered_10b[1239] = 10'h3F0;
    I_filtered_10b[1238] = 10'h3E9;
    I_filtered_10b[1237] = 10'h3E0;
    I_filtered_10b[1236] = 10'h3DC;
    I_filtered_10b[1235] = 10'h3D7;
    I_filtered_10b[1234] = 10'h3D8;
    I_filtered_10b[1233] = 10'h3D7;
    I_filtered_10b[1232] = 10'h3DB;
    I_filtered_10b[1231] = 10'h3E0;
    I_filtered_10b[1230] = 10'h3E7;
    I_filtered_10b[1229] = 10'h3EE;
    I_filtered_10b[1228] = 10'h3F2;
    I_filtered_10b[1227] = 10'h3F9;
    I_filtered_10b[1226] = 10'h3FC;
    I_filtered_10b[1225] = 10'h000;
    I_filtered_10b[1224] = 10'h000;
    I_filtered_10b[1223] = 10'h000;
    I_filtered_10b[1222] = 10'h001;
    I_filtered_10b[1221] = 10'h003;
    I_filtered_10b[1220] = 10'h004;
    I_filtered_10b[1219] = 10'h009;
    I_filtered_10b[1218] = 10'h00E;
    I_filtered_10b[1217] = 10'h015;
    I_filtered_10b[1216] = 10'h022;
    I_filtered_10b[1215] = 10'h02E;
    I_filtered_10b[1214] = 10'h03E;
    I_filtered_10b[1213] = 10'h050;
    I_filtered_10b[1212] = 10'h066;
    I_filtered_10b[1211] = 10'h07A;
    I_filtered_10b[1210] = 10'h08F;
    I_filtered_10b[1209] = 10'h0A2;
    I_filtered_10b[1208] = 10'h0B2;
    I_filtered_10b[1207] = 10'h0BF;
    I_filtered_10b[1206] = 10'h0C8;
    I_filtered_10b[1205] = 10'h0CC;
    I_filtered_10b[1204] = 10'h0CC;
    I_filtered_10b[1203] = 10'h0CA;
    I_filtered_10b[1202] = 10'h0C4;
    I_filtered_10b[1201] = 10'h0BC;
    I_filtered_10b[1200] = 10'h0B4;
    I_filtered_10b[1199] = 10'h0AA;
    I_filtered_10b[1198] = 10'h0A1;
    I_filtered_10b[1197] = 10'h09B;
    I_filtered_10b[1196] = 10'h095;
    I_filtered_10b[1195] = 10'h094;
    I_filtered_10b[1194] = 10'h092;
    I_filtered_10b[1193] = 10'h08E;
    I_filtered_10b[1192] = 10'h08D;
    I_filtered_10b[1191] = 10'h08B;
    I_filtered_10b[1190] = 10'h083;
    I_filtered_10b[1189] = 10'h078;
    I_filtered_10b[1188] = 10'h06A;
    I_filtered_10b[1187] = 10'h057;
    I_filtered_10b[1186] = 10'h040;
    I_filtered_10b[1185] = 10'h027;
    I_filtered_10b[1184] = 10'h00C;
    I_filtered_10b[1183] = 10'h3F2;
    I_filtered_10b[1182] = 10'h3DD;
    I_filtered_10b[1181] = 10'h3CC;
    I_filtered_10b[1180] = 10'h3C1;
    I_filtered_10b[1179] = 10'h3BC;
    I_filtered_10b[1178] = 10'h3C2;
    I_filtered_10b[1177] = 10'h3CF;
    I_filtered_10b[1176] = 10'h3E4;
    I_filtered_10b[1175] = 10'h3FC;
    I_filtered_10b[1174] = 10'h01C;
    I_filtered_10b[1173] = 10'h03F;
    I_filtered_10b[1172] = 10'h060;
    I_filtered_10b[1171] = 10'h081;
    I_filtered_10b[1170] = 10'h09C;
    I_filtered_10b[1169] = 10'h0B2;
    I_filtered_10b[1168] = 10'h0C4;
    I_filtered_10b[1167] = 10'h0CF;
    I_filtered_10b[1166] = 10'h0D2;
    I_filtered_10b[1165] = 10'h0D2;
    I_filtered_10b[1164] = 10'h0CF;
    I_filtered_10b[1163] = 10'h0C8;
    I_filtered_10b[1162] = 10'h0BD;
    I_filtered_10b[1161] = 10'h0B5;
    I_filtered_10b[1160] = 10'h0A9;
    I_filtered_10b[1159] = 10'h0A0;
    I_filtered_10b[1158] = 10'h09A;
    I_filtered_10b[1157] = 10'h092;
    I_filtered_10b[1156] = 10'h08F;
    I_filtered_10b[1155] = 10'h08C;
    I_filtered_10b[1154] = 10'h088;
    I_filtered_10b[1153] = 10'h087;
    I_filtered_10b[1152] = 10'h085;
    I_filtered_10b[1151] = 10'h080;
    I_filtered_10b[1150] = 10'h079;
    I_filtered_10b[1149] = 10'h071;
    I_filtered_10b[1148] = 10'h066;
    I_filtered_10b[1147] = 10'h058;
    I_filtered_10b[1146] = 10'h04A;
    I_filtered_10b[1145] = 10'h039;
    I_filtered_10b[1144] = 10'h02A;
    I_filtered_10b[1143] = 10'h01E;
    I_filtered_10b[1142] = 10'h014;
    I_filtered_10b[1141] = 10'h00C;
    I_filtered_10b[1140] = 10'h008;
    I_filtered_10b[1139] = 10'h009;
    I_filtered_10b[1138] = 10'h00C;
    I_filtered_10b[1137] = 10'h013;
    I_filtered_10b[1136] = 10'h01A;
    I_filtered_10b[1135] = 10'h025;
    I_filtered_10b[1134] = 10'h030;
    I_filtered_10b[1133] = 10'h03B;
    I_filtered_10b[1132] = 10'h043;
    I_filtered_10b[1131] = 10'h04A;
    I_filtered_10b[1130] = 10'h04C;
    I_filtered_10b[1129] = 10'h04F;
    I_filtered_10b[1128] = 10'h04F;
    I_filtered_10b[1127] = 10'h04D;
    I_filtered_10b[1126] = 10'h04B;
    I_filtered_10b[1125] = 10'h04D;
    I_filtered_10b[1124] = 10'h051;
    I_filtered_10b[1123] = 10'h055;
    I_filtered_10b[1122] = 10'h05E;
    I_filtered_10b[1121] = 10'h067;
    I_filtered_10b[1120] = 10'h074;
    I_filtered_10b[1119] = 10'h082;
    I_filtered_10b[1118] = 10'h08E;
    I_filtered_10b[1117] = 10'h09A;
    I_filtered_10b[1116] = 10'h0A3;
    I_filtered_10b[1115] = 10'h0A5;
    I_filtered_10b[1114] = 10'h0A5;
    I_filtered_10b[1113] = 10'h09F;
    I_filtered_10b[1112] = 10'h08F;
    I_filtered_10b[1111] = 10'h079;
    I_filtered_10b[1110] = 10'h05D;
    I_filtered_10b[1109] = 10'h03A;
    I_filtered_10b[1108] = 10'h011;
    I_filtered_10b[1107] = 10'h3E8;
    I_filtered_10b[1106] = 10'h3BD;
    I_filtered_10b[1105] = 10'h396;
    I_filtered_10b[1104] = 10'h377;
    I_filtered_10b[1103] = 10'h35E;
    I_filtered_10b[1102] = 10'h34F;
    I_filtered_10b[1101] = 10'h349;
    I_filtered_10b[1100] = 10'h350;
    I_filtered_10b[1099] = 10'h35D;
    I_filtered_10b[1098] = 10'h373;
    I_filtered_10b[1097] = 10'h38F;
    I_filtered_10b[1096] = 10'h3AF;
    I_filtered_10b[1095] = 10'h3D1;
    I_filtered_10b[1094] = 10'h3F0;
    I_filtered_10b[1093] = 10'h00D;
    I_filtered_10b[1092] = 10'h025;
    I_filtered_10b[1091] = 10'h038;
    I_filtered_10b[1090] = 10'h047;
    I_filtered_10b[1089] = 10'h054;
    I_filtered_10b[1088] = 10'h059;
    I_filtered_10b[1087] = 10'h05E;
    I_filtered_10b[1086] = 10'h066;
    I_filtered_10b[1085] = 10'h06B;
    I_filtered_10b[1084] = 10'h070;
    I_filtered_10b[1083] = 10'h07A;
    I_filtered_10b[1082] = 10'h085;
    I_filtered_10b[1081] = 10'h090;
    I_filtered_10b[1080] = 10'h0A0;
    I_filtered_10b[1079] = 10'h0AC;
    I_filtered_10b[1078] = 10'h0B8;
    I_filtered_10b[1077] = 10'h0C2;
    I_filtered_10b[1076] = 10'h0C8;
    I_filtered_10b[1075] = 10'h0CC;
    I_filtered_10b[1074] = 10'h0CB;
    I_filtered_10b[1073] = 10'h0C7;
    I_filtered_10b[1072] = 10'h0BD;
    I_filtered_10b[1071] = 10'h0B2;
    I_filtered_10b[1070] = 10'h0A4;
    I_filtered_10b[1069] = 10'h096;
    I_filtered_10b[1068] = 10'h08A;
    I_filtered_10b[1067] = 10'h07B;
    I_filtered_10b[1066] = 10'h071;
    I_filtered_10b[1065] = 10'h066;
    I_filtered_10b[1064] = 10'h05F;
    I_filtered_10b[1063] = 10'h054;
    I_filtered_10b[1062] = 10'h04D;
    I_filtered_10b[1061] = 10'h045;
    I_filtered_10b[1060] = 10'h03C;
    I_filtered_10b[1059] = 10'h036;
    I_filtered_10b[1058] = 10'h02E;
    I_filtered_10b[1057] = 10'h027;
    I_filtered_10b[1056] = 10'h01E;
    I_filtered_10b[1055] = 10'h01A;
    I_filtered_10b[1054] = 10'h011;
    I_filtered_10b[1053] = 10'h00B;
    I_filtered_10b[1052] = 10'h004;
    I_filtered_10b[1051] = 10'h3FE;
    I_filtered_10b[1050] = 10'h3F5;
    I_filtered_10b[1049] = 10'h3EC;
    I_filtered_10b[1048] = 10'h3E4;
    I_filtered_10b[1047] = 10'h3D6;
    I_filtered_10b[1046] = 10'h3CB;
    I_filtered_10b[1045] = 10'h3BB;
    I_filtered_10b[1044] = 10'h3AB;
    I_filtered_10b[1043] = 10'h398;
    I_filtered_10b[1042] = 10'h388;
    I_filtered_10b[1041] = 10'h373;
    I_filtered_10b[1040] = 10'h361;
    I_filtered_10b[1039] = 10'h34E;
    I_filtered_10b[1038] = 10'h340;
    I_filtered_10b[1037] = 10'h335;
    I_filtered_10b[1036] = 10'h32E;
    I_filtered_10b[1035] = 10'h32B;
    I_filtered_10b[1034] = 10'h32E;
    I_filtered_10b[1033] = 10'h338;
    I_filtered_10b[1032] = 10'h345;
    I_filtered_10b[1031] = 10'h357;
    I_filtered_10b[1030] = 10'h368;
    I_filtered_10b[1029] = 10'h37B;
    I_filtered_10b[1028] = 10'h390;
    I_filtered_10b[1027] = 10'h3A1;
    I_filtered_10b[1026] = 10'h3B1;
    I_filtered_10b[1025] = 10'h3BD;
    I_filtered_10b[1024] = 10'h3C7;
    I_filtered_10b[1023] = 10'h3CB;
    I_filtered_10b[1022] = 10'h3CD;
    I_filtered_10b[1021] = 10'h3C7;
    I_filtered_10b[1020] = 10'h3BB;
    I_filtered_10b[1019] = 10'h3AD;
    I_filtered_10b[1018] = 10'h398;
    I_filtered_10b[1017] = 10'h383;
    I_filtered_10b[1016] = 10'h369;
    I_filtered_10b[1015] = 10'h350;
    I_filtered_10b[1014] = 10'h33A;
    I_filtered_10b[1013] = 10'h325;
    I_filtered_10b[1012] = 10'h317;
    I_filtered_10b[1011] = 10'h313;
    I_filtered_10b[1010] = 10'h316;
    I_filtered_10b[1009] = 10'h320;
    I_filtered_10b[1008] = 10'h337;
    I_filtered_10b[1007] = 10'h357;
    I_filtered_10b[1006] = 10'h381;
    I_filtered_10b[1005] = 10'h3B0;
    I_filtered_10b[1004] = 10'h3E7;
    I_filtered_10b[1003] = 10'h01C;
    I_filtered_10b[1002] = 10'h055;
    I_filtered_10b[1001] = 10'h088;
    I_filtered_10b[1000] = 10'h0B6;
    I_filtered_10b[999] = 10'h0D9;
    I_filtered_10b[998] = 10'h0F1;
    I_filtered_10b[997] = 10'h0FC;
    I_filtered_10b[996] = 10'h0FB;
    I_filtered_10b[995] = 10'h0EE;
    I_filtered_10b[994] = 10'h0D2;
    I_filtered_10b[993] = 10'h0AE;
    I_filtered_10b[992] = 10'h082;
    I_filtered_10b[991] = 10'h053;
    I_filtered_10b[990] = 10'h022;
    I_filtered_10b[989] = 10'h3F3;
    I_filtered_10b[988] = 10'h3CB;
    I_filtered_10b[987] = 10'h3A9;
    I_filtered_10b[986] = 10'h38F;
    I_filtered_10b[985] = 10'h380;
    I_filtered_10b[984] = 10'h37D;
    I_filtered_10b[983] = 10'h381;
    I_filtered_10b[982] = 10'h38F;
    I_filtered_10b[981] = 10'h3A5;
    I_filtered_10b[980] = 10'h3C4;
    I_filtered_10b[979] = 10'h3E5;
    I_filtered_10b[978] = 10'h00C;
    I_filtered_10b[977] = 10'h032;
    I_filtered_10b[976] = 10'h056;
    I_filtered_10b[975] = 10'h078;
    I_filtered_10b[974] = 10'h092;
    I_filtered_10b[973] = 10'h0A7;
    I_filtered_10b[972] = 10'h0B1;
    I_filtered_10b[971] = 10'h0B1;
    I_filtered_10b[970] = 10'h0A9;
    I_filtered_10b[969] = 10'h09A;
    I_filtered_10b[968] = 10'h085;
    I_filtered_10b[967] = 10'h069;
    I_filtered_10b[966] = 10'h04C;
    I_filtered_10b[965] = 10'h02A;
    I_filtered_10b[964] = 10'h00D;
    I_filtered_10b[963] = 10'h3F0;
    I_filtered_10b[962] = 10'h3D6;
    I_filtered_10b[961] = 10'h3C0;
    I_filtered_10b[960] = 10'h3AE;
    I_filtered_10b[959] = 10'h3A1;
    I_filtered_10b[958] = 10'h39B;
    I_filtered_10b[957] = 10'h397;
    I_filtered_10b[956] = 10'h396;
    I_filtered_10b[955] = 10'h399;
    I_filtered_10b[954] = 10'h39F;
    I_filtered_10b[953] = 10'h3A4;
    I_filtered_10b[952] = 10'h3A9;
    I_filtered_10b[951] = 10'h3AF;
    I_filtered_10b[950] = 10'h3B3;
    I_filtered_10b[949] = 10'h3B6;
    I_filtered_10b[948] = 10'h3B9;
    I_filtered_10b[947] = 10'h3BB;
    I_filtered_10b[946] = 10'h3BB;
    I_filtered_10b[945] = 10'h3B9;
    I_filtered_10b[944] = 10'h3B8;
    I_filtered_10b[943] = 10'h3B3;
    I_filtered_10b[942] = 10'h3AE;
    I_filtered_10b[941] = 10'h3A6;
    I_filtered_10b[940] = 10'h39E;
    I_filtered_10b[939] = 10'h395;
    I_filtered_10b[938] = 10'h38B;
    I_filtered_10b[937] = 10'h380;
    I_filtered_10b[936] = 10'h376;
    I_filtered_10b[935] = 10'h36B;
    I_filtered_10b[934] = 10'h363;
    I_filtered_10b[933] = 10'h361;
    I_filtered_10b[932] = 10'h361;
    I_filtered_10b[931] = 10'h365;
    I_filtered_10b[930] = 10'h371;
    I_filtered_10b[929] = 10'h383;
    I_filtered_10b[928] = 10'h39A;
    I_filtered_10b[927] = 10'h3B6;
    I_filtered_10b[926] = 10'h3D6;
    I_filtered_10b[925] = 10'h3F7;
    I_filtered_10b[924] = 10'h01A;
    I_filtered_10b[923] = 10'h03A;
    I_filtered_10b[922] = 10'h055;
    I_filtered_10b[921] = 10'h06A;
    I_filtered_10b[920] = 10'h078;
    I_filtered_10b[919] = 10'h07D;
    I_filtered_10b[918] = 10'h079;
    I_filtered_10b[917] = 10'h06D;
    I_filtered_10b[916] = 10'h057;
    I_filtered_10b[915] = 10'h03D;
    I_filtered_10b[914] = 10'h01C;
    I_filtered_10b[913] = 10'h3F9;
    I_filtered_10b[912] = 10'h3D7;
    I_filtered_10b[911] = 10'h3B4;
    I_filtered_10b[910] = 10'h398;
    I_filtered_10b[909] = 10'h37F;
    I_filtered_10b[908] = 10'h36C;
    I_filtered_10b[907] = 10'h35F;
    I_filtered_10b[906] = 10'h35B;
    I_filtered_10b[905] = 10'h35B;
    I_filtered_10b[904] = 10'h361;
    I_filtered_10b[903] = 10'h36D;
    I_filtered_10b[902] = 10'h37E;
    I_filtered_10b[901] = 10'h38F;
    I_filtered_10b[900] = 10'h3A2;
    I_filtered_10b[899] = 10'h3B5;
    I_filtered_10b[898] = 10'h3C8;
    I_filtered_10b[897] = 10'h3D9;
    I_filtered_10b[896] = 10'h3E9;
    I_filtered_10b[895] = 10'h3F4;
    I_filtered_10b[894] = 10'h3FC;
    I_filtered_10b[893] = 10'h3FE;
    I_filtered_10b[892] = 10'h3FF;
    I_filtered_10b[891] = 10'h3F9;
    I_filtered_10b[890] = 10'h3EE;
    I_filtered_10b[889] = 10'h3DF;
    I_filtered_10b[888] = 10'h3CC;
    I_filtered_10b[887] = 10'h3B5;
    I_filtered_10b[886] = 10'h39B;
    I_filtered_10b[885] = 10'h384;
    I_filtered_10b[884] = 10'h36D;
    I_filtered_10b[883] = 10'h35C;
    I_filtered_10b[882] = 10'h34E;
    I_filtered_10b[881] = 10'h34B;
    I_filtered_10b[880] = 10'h34F;
    I_filtered_10b[879] = 10'h35C;
    I_filtered_10b[878] = 10'h373;
    I_filtered_10b[877] = 10'h38F;
    I_filtered_10b[876] = 10'h3B3;
    I_filtered_10b[875] = 10'h3DA;
    I_filtered_10b[874] = 10'h007;
    I_filtered_10b[873] = 10'h02F;
    I_filtered_10b[872] = 10'h05A;
    I_filtered_10b[871] = 10'h07F;
    I_filtered_10b[870] = 10'h09F;
    I_filtered_10b[869] = 10'h0B9;
    I_filtered_10b[868] = 10'h0CD;
    I_filtered_10b[867] = 10'h0D8;
    I_filtered_10b[866] = 10'h0DE;
    I_filtered_10b[865] = 10'h0E1;
    I_filtered_10b[864] = 10'h0DD;
    I_filtered_10b[863] = 10'h0D6;
    I_filtered_10b[862] = 10'h0CF;
    I_filtered_10b[861] = 10'h0CA;
    I_filtered_10b[860] = 10'h0C4;
    I_filtered_10b[859] = 10'h0C0;
    I_filtered_10b[858] = 10'h0BF;
    I_filtered_10b[857] = 10'h0BD;
    I_filtered_10b[856] = 10'h0BC;
    I_filtered_10b[855] = 10'h0BA;
    I_filtered_10b[854] = 10'h0BA;
    I_filtered_10b[853] = 10'h0B6;
    I_filtered_10b[852] = 10'h0B4;
    I_filtered_10b[851] = 10'h0B1;
    I_filtered_10b[850] = 10'h0AF;
    I_filtered_10b[849] = 10'h0AC;
    I_filtered_10b[848] = 10'h0A9;
    I_filtered_10b[847] = 10'h0AA;
    I_filtered_10b[846] = 10'h0A9;
    I_filtered_10b[845] = 10'h0AA;
    I_filtered_10b[844] = 10'h0AC;
    I_filtered_10b[843] = 10'h0AD;
    I_filtered_10b[842] = 10'h0A6;
    I_filtered_10b[841] = 10'h09F;
    I_filtered_10b[840] = 10'h094;
    I_filtered_10b[839] = 10'h07F;
    I_filtered_10b[838] = 10'h066;
    I_filtered_10b[837] = 10'h046;
    I_filtered_10b[836] = 10'h021;
    I_filtered_10b[835] = 10'h3F4;
    I_filtered_10b[834] = 10'h3C8;
    I_filtered_10b[833] = 10'h399;
    I_filtered_10b[832] = 10'h36D;
    I_filtered_10b[831] = 10'h349;
    I_filtered_10b[830] = 10'h32C;
    I_filtered_10b[829] = 10'h319;
    I_filtered_10b[828] = 10'h310;
    I_filtered_10b[827] = 10'h315;
    I_filtered_10b[826] = 10'h321;
    I_filtered_10b[825] = 10'h337;
    I_filtered_10b[824] = 10'h353;
    I_filtered_10b[823] = 10'h374;
    I_filtered_10b[822] = 10'h398;
    I_filtered_10b[821] = 10'h3B8;
    I_filtered_10b[820] = 10'h3D6;
    I_filtered_10b[819] = 10'h3EE;
    I_filtered_10b[818] = 10'h3FF;
    I_filtered_10b[817] = 10'h00E;
    I_filtered_10b[816] = 10'h01A;
    I_filtered_10b[815] = 10'h020;
    I_filtered_10b[814] = 10'h025;
    I_filtered_10b[813] = 10'h02F;
    I_filtered_10b[812] = 10'h039;
    I_filtered_10b[811] = 10'h042;
    I_filtered_10b[810] = 10'h053;
    I_filtered_10b[809] = 10'h066;
    I_filtered_10b[808] = 10'h07A;
    I_filtered_10b[807] = 10'h092;
    I_filtered_10b[806] = 10'h0A7;
    I_filtered_10b[805] = 10'h0BA;
    I_filtered_10b[804] = 10'h0C9;
    I_filtered_10b[803] = 10'h0D2;
    I_filtered_10b[802] = 10'h0D8;
    I_filtered_10b[801] = 10'h0D5;
    I_filtered_10b[800] = 10'h0CE;
    I_filtered_10b[799] = 10'h0BF;
    I_filtered_10b[798] = 10'h0AD;
    I_filtered_10b[797] = 10'h096;
    I_filtered_10b[796] = 10'h080;
    I_filtered_10b[795] = 10'h06B;
    I_filtered_10b[794] = 10'h054;
    I_filtered_10b[793] = 10'h043;
    I_filtered_10b[792] = 10'h034;
    I_filtered_10b[791] = 10'h028;
    I_filtered_10b[790] = 10'h01B;
    I_filtered_10b[789] = 10'h014;
    I_filtered_10b[788] = 10'h00B;
    I_filtered_10b[787] = 10'h003;
    I_filtered_10b[786] = 10'h3FD;
    I_filtered_10b[785] = 10'h3F7;
    I_filtered_10b[784] = 10'h3F0;
    I_filtered_10b[783] = 10'h3E7;
    I_filtered_10b[782] = 10'h3E2;
    I_filtered_10b[781] = 10'h3D8;
    I_filtered_10b[780] = 10'h3D1;
    I_filtered_10b[779] = 10'h3C9;
    I_filtered_10b[778] = 10'h3C3;
    I_filtered_10b[777] = 10'h3BB;
    I_filtered_10b[776] = 10'h3B3;
    I_filtered_10b[775] = 10'h3AD;
    I_filtered_10b[774] = 10'h3A3;
    I_filtered_10b[773] = 10'h39B;
    I_filtered_10b[772] = 10'h391;
    I_filtered_10b[771] = 10'h386;
    I_filtered_10b[770] = 10'h378;
    I_filtered_10b[769] = 10'h36C;
    I_filtered_10b[768] = 10'h35D;
    I_filtered_10b[767] = 10'h34E;
    I_filtered_10b[766] = 10'h340;
    I_filtered_10b[765] = 10'h336;
    I_filtered_10b[764] = 10'h330;
    I_filtered_10b[763] = 10'h32E;
    I_filtered_10b[762] = 10'h331;
    I_filtered_10b[761] = 10'h339;
    I_filtered_10b[760] = 10'h347;
    I_filtered_10b[759] = 10'h358;
    I_filtered_10b[758] = 10'h36D;
    I_filtered_10b[757] = 10'h386;
    I_filtered_10b[756] = 10'h39E;
    I_filtered_10b[755] = 10'h3B6;
    I_filtered_10b[754] = 10'h3CC;
    I_filtered_10b[753] = 10'h3DC;
    I_filtered_10b[752] = 10'h3E9;
    I_filtered_10b[751] = 10'h3F4;
    I_filtered_10b[750] = 10'h3F8;
    I_filtered_10b[749] = 10'h3F8;
    I_filtered_10b[748] = 10'h3F7;
    I_filtered_10b[747] = 10'h3F4;
    I_filtered_10b[746] = 10'h3F0;
    I_filtered_10b[745] = 10'h3EC;
    I_filtered_10b[744] = 10'h3E7;
    I_filtered_10b[743] = 10'h3E4;
    I_filtered_10b[742] = 10'h3E5;
    I_filtered_10b[741] = 10'h3E6;
    I_filtered_10b[740] = 10'h3EA;
    I_filtered_10b[739] = 10'h3EC;
    I_filtered_10b[738] = 10'h3EF;
    I_filtered_10b[737] = 10'h3F2;
    I_filtered_10b[736] = 10'h3F3;
    I_filtered_10b[735] = 10'h3EE;
    I_filtered_10b[734] = 10'h3E5;
    I_filtered_10b[733] = 10'h3DB;
    I_filtered_10b[732] = 10'h3CA;
    I_filtered_10b[731] = 10'h3B9;
    I_filtered_10b[730] = 10'h3A5;
    I_filtered_10b[729] = 10'h38F;
    I_filtered_10b[728] = 10'h37E;
    I_filtered_10b[727] = 10'h36E;
    I_filtered_10b[726] = 10'h362;
    I_filtered_10b[725] = 10'h35C;
    I_filtered_10b[724] = 10'h35B;
    I_filtered_10b[723] = 10'h360;
    I_filtered_10b[722] = 10'h36D;
    I_filtered_10b[721] = 10'h380;
    I_filtered_10b[720] = 10'h398;
    I_filtered_10b[719] = 10'h3B4;
    I_filtered_10b[718] = 10'h3D6;
    I_filtered_10b[717] = 10'h3F7;
    I_filtered_10b[716] = 10'h018;
    I_filtered_10b[715] = 10'h036;
    I_filtered_10b[714] = 10'h04D;
    I_filtered_10b[713] = 10'h061;
    I_filtered_10b[712] = 10'h06D;
    I_filtered_10b[711] = 10'h071;
    I_filtered_10b[710] = 10'h06E;
    I_filtered_10b[709] = 10'h067;
    I_filtered_10b[708] = 10'h05A;
    I_filtered_10b[707] = 10'h04A;
    I_filtered_10b[706] = 10'h039;
    I_filtered_10b[705] = 10'h026;
    I_filtered_10b[704] = 10'h016;
    I_filtered_10b[703] = 10'h008;
    I_filtered_10b[702] = 10'h3FD;
    I_filtered_10b[701] = 10'h3F5;
    I_filtered_10b[700] = 10'h3EE;
    I_filtered_10b[699] = 10'h3E8;
    I_filtered_10b[698] = 10'h3E6;
    I_filtered_10b[697] = 10'h3E3;
    I_filtered_10b[696] = 10'h3DD;
    I_filtered_10b[695] = 10'h3D6;
    I_filtered_10b[694] = 10'h3CF;
    I_filtered_10b[693] = 10'h3C2;
    I_filtered_10b[692] = 10'h3B6;
    I_filtered_10b[691] = 10'h3A8;
    I_filtered_10b[690] = 10'h397;
    I_filtered_10b[689] = 10'h38A;
    I_filtered_10b[688] = 10'h37D;
    I_filtered_10b[687] = 10'h373;
    I_filtered_10b[686] = 10'h36C;
    I_filtered_10b[685] = 10'h367;
    I_filtered_10b[684] = 10'h367;
    I_filtered_10b[683] = 10'h36B;
    I_filtered_10b[682] = 10'h375;
    I_filtered_10b[681] = 10'h381;
    I_filtered_10b[680] = 10'h391;
    I_filtered_10b[679] = 10'h3A2;
    I_filtered_10b[678] = 10'h3B4;
    I_filtered_10b[677] = 10'h3C7;
    I_filtered_10b[676] = 10'h3D6;
    I_filtered_10b[675] = 10'h3E3;
    I_filtered_10b[674] = 10'h3ED;
    I_filtered_10b[673] = 10'h3F5;
    I_filtered_10b[672] = 10'h3F8;
    I_filtered_10b[671] = 10'h3F9;
    I_filtered_10b[670] = 10'h3F5;
    I_filtered_10b[669] = 10'h3EF;
    I_filtered_10b[668] = 10'h3E6;
    I_filtered_10b[667] = 10'h3DB;
    I_filtered_10b[666] = 10'h3CF;
    I_filtered_10b[665] = 10'h3C2;
    I_filtered_10b[664] = 10'h3B7;
    I_filtered_10b[663] = 10'h3AD;
    I_filtered_10b[662] = 10'h3A6;
    I_filtered_10b[661] = 10'h3A0;
    I_filtered_10b[660] = 10'h39F;
    I_filtered_10b[659] = 10'h3A1;
    I_filtered_10b[658] = 10'h3A5;
    I_filtered_10b[657] = 10'h3AD;
    I_filtered_10b[656] = 10'h3B6;
    I_filtered_10b[655] = 10'h3C3;
    I_filtered_10b[654] = 10'h3D0;
    I_filtered_10b[653] = 10'h3E1;
    I_filtered_10b[652] = 10'h3EF;
    I_filtered_10b[651] = 10'h3FD;
    I_filtered_10b[650] = 10'h00B;
    I_filtered_10b[649] = 10'h015;
    I_filtered_10b[648] = 10'h01E;
    I_filtered_10b[647] = 10'h023;
    I_filtered_10b[646] = 10'h026;
    I_filtered_10b[645] = 10'h024;
    I_filtered_10b[644] = 10'h024;
    I_filtered_10b[643] = 10'h022;
    I_filtered_10b[642] = 10'h01F;
    I_filtered_10b[641] = 10'h01E;
    I_filtered_10b[640] = 10'h01C;
    I_filtered_10b[639] = 10'h01D;
    I_filtered_10b[638] = 10'h020;
    I_filtered_10b[637] = 10'h023;
    I_filtered_10b[636] = 10'h028;
    I_filtered_10b[635] = 10'h02B;
    I_filtered_10b[634] = 10'h02B;
    I_filtered_10b[633] = 10'h02C;
    I_filtered_10b[632] = 10'h028;
    I_filtered_10b[631] = 10'h01F;
    I_filtered_10b[630] = 10'h012;
    I_filtered_10b[629] = 10'h002;
    I_filtered_10b[628] = 10'h3ED;
    I_filtered_10b[627] = 10'h3D4;
    I_filtered_10b[626] = 10'h3B9;
    I_filtered_10b[625] = 10'h39F;
    I_filtered_10b[624] = 10'h386;
    I_filtered_10b[623] = 10'h374;
    I_filtered_10b[622] = 10'h365;
    I_filtered_10b[621] = 10'h35D;
    I_filtered_10b[620] = 10'h35B;
    I_filtered_10b[619] = 10'h362;
    I_filtered_10b[618] = 10'h36C;
    I_filtered_10b[617] = 10'h37C;
    I_filtered_10b[616] = 10'h38F;
    I_filtered_10b[615] = 10'h3A5;
    I_filtered_10b[614] = 10'h3BD;
    I_filtered_10b[613] = 10'h3D1;
    I_filtered_10b[612] = 10'h3E5;
    I_filtered_10b[611] = 10'h3F5;
    I_filtered_10b[610] = 10'h000;
    I_filtered_10b[609] = 10'h00B;
    I_filtered_10b[608] = 10'h014;
    I_filtered_10b[607] = 10'h01A;
    I_filtered_10b[606] = 10'h01F;
    I_filtered_10b[605] = 10'h029;
    I_filtered_10b[604] = 10'h034;
    I_filtered_10b[603] = 10'h040;
    I_filtered_10b[602] = 10'h051;
    I_filtered_10b[601] = 10'h064;
    I_filtered_10b[600] = 10'h077;
    I_filtered_10b[599] = 10'h091;
    I_filtered_10b[598] = 10'h0A5;
    I_filtered_10b[597] = 10'h0BC;
    I_filtered_10b[596] = 10'h0CC;
    I_filtered_10b[595] = 10'h0D7;
    I_filtered_10b[594] = 10'h0DE;
    I_filtered_10b[593] = 10'h0DE;
    I_filtered_10b[592] = 10'h0D5;
    I_filtered_10b[591] = 10'h0C2;
    I_filtered_10b[590] = 10'h0AA;
    I_filtered_10b[589] = 10'h08A;
    I_filtered_10b[588] = 10'h069;
    I_filtered_10b[587] = 10'h045;
    I_filtered_10b[586] = 10'h01F;
    I_filtered_10b[585] = 10'h000;
    I_filtered_10b[584] = 10'h3E2;
    I_filtered_10b[583] = 10'h3CC;
    I_filtered_10b[582] = 10'h3BD;
    I_filtered_10b[581] = 10'h3B6;
    I_filtered_10b[580] = 10'h3B7;
    I_filtered_10b[579] = 10'h3C2;
    I_filtered_10b[578] = 10'h3D8;
    I_filtered_10b[577] = 10'h3F4;
    I_filtered_10b[576] = 10'h017;
    I_filtered_10b[575] = 10'h03D;
    I_filtered_10b[574] = 10'h067;
    I_filtered_10b[573] = 10'h090;
    I_filtered_10b[572] = 10'h0B4;
    I_filtered_10b[571] = 10'h0D4;
    I_filtered_10b[570] = 10'h0EB;
    I_filtered_10b[569] = 10'h0F6;
    I_filtered_10b[568] = 10'h0F6;
    I_filtered_10b[567] = 10'h0ED;
    I_filtered_10b[566] = 10'h0D6;
    I_filtered_10b[565] = 10'h0B4;
    I_filtered_10b[564] = 10'h087;
    I_filtered_10b[563] = 10'h055;
    I_filtered_10b[562] = 10'h019;
    I_filtered_10b[561] = 10'h3E0;
    I_filtered_10b[560] = 10'h3A6;
    I_filtered_10b[559] = 10'h370;
    I_filtered_10b[558] = 10'h344;
    I_filtered_10b[557] = 10'h321;
    I_filtered_10b[556] = 10'h30B;
    I_filtered_10b[555] = 10'h304;
    I_filtered_10b[554] = 10'h309;
    I_filtered_10b[553] = 10'h319;
    I_filtered_10b[552] = 10'h335;
    I_filtered_10b[551] = 10'h359;
    I_filtered_10b[550] = 10'h383;
    I_filtered_10b[549] = 10'h3B2;
    I_filtered_10b[548] = 10'h3DE;
    I_filtered_10b[547] = 10'h007;
    I_filtered_10b[546] = 10'h02C;
    I_filtered_10b[545] = 10'h048;
    I_filtered_10b[544] = 10'h05F;
    I_filtered_10b[543] = 10'h06E;
    I_filtered_10b[542] = 10'h071;
    I_filtered_10b[541] = 10'h070;
    I_filtered_10b[540] = 10'h06B;
    I_filtered_10b[539] = 10'h062;
    I_filtered_10b[538] = 10'h054;
    I_filtered_10b[537] = 10'h049;
    I_filtered_10b[536] = 10'h03D;
    I_filtered_10b[535] = 10'h033;
    I_filtered_10b[534] = 10'h02C;
    I_filtered_10b[533] = 10'h026;
    I_filtered_10b[532] = 10'h020;
    I_filtered_10b[531] = 10'h01D;
    I_filtered_10b[530] = 10'h019;
    I_filtered_10b[529] = 10'h01A;
    I_filtered_10b[528] = 10'h017;
    I_filtered_10b[527] = 10'h014;
    I_filtered_10b[526] = 10'h011;
    I_filtered_10b[525] = 10'h00F;
    I_filtered_10b[524] = 10'h009;
    I_filtered_10b[523] = 10'h004;
    I_filtered_10b[522] = 10'h000;
    I_filtered_10b[521] = 10'h3FB;
    I_filtered_10b[520] = 10'h3F8;
    I_filtered_10b[519] = 10'h3F6;
    I_filtered_10b[518] = 10'h3F4;
    I_filtered_10b[517] = 10'h3F0;
    I_filtered_10b[516] = 10'h3EC;
    I_filtered_10b[515] = 10'h3E9;
    I_filtered_10b[514] = 10'h3E1;
    I_filtered_10b[513] = 10'h3D9;
    I_filtered_10b[512] = 10'h3CE;
    I_filtered_10b[511] = 10'h3C2;
    I_filtered_10b[510] = 10'h3B4;
    I_filtered_10b[509] = 10'h3A6;
    I_filtered_10b[508] = 10'h395;
    I_filtered_10b[507] = 10'h386;
    I_filtered_10b[506] = 10'h377;
    I_filtered_10b[505] = 10'h36C;
    I_filtered_10b[504] = 10'h365;
    I_filtered_10b[503] = 10'h361;
    I_filtered_10b[502] = 10'h362;
    I_filtered_10b[501] = 10'h36A;
    I_filtered_10b[500] = 10'h378;
    I_filtered_10b[499] = 10'h38A;
    I_filtered_10b[498] = 10'h3A1;
    I_filtered_10b[497] = 10'h3BA;
    I_filtered_10b[496] = 10'h3D4;
    I_filtered_10b[495] = 10'h3F0;
    I_filtered_10b[494] = 10'h007;
    I_filtered_10b[493] = 10'h01D;
    I_filtered_10b[492] = 10'h02D;
    I_filtered_10b[491] = 10'h039;
    I_filtered_10b[490] = 10'h03E;
    I_filtered_10b[489] = 10'h03D;
    I_filtered_10b[488] = 10'h035;
    I_filtered_10b[487] = 10'h024;
    I_filtered_10b[486] = 10'h010;
    I_filtered_10b[485] = 10'h3F6;
    I_filtered_10b[484] = 10'h3D7;
    I_filtered_10b[483] = 10'h3B5;
    I_filtered_10b[482] = 10'h397;
    I_filtered_10b[481] = 10'h37A;
    I_filtered_10b[480] = 10'h365;
    I_filtered_10b[479] = 10'h353;
    I_filtered_10b[478] = 10'h34D;
    I_filtered_10b[477] = 10'h34F;
    I_filtered_10b[476] = 10'h35A;
    I_filtered_10b[475] = 10'h36D;
    I_filtered_10b[474] = 10'h386;
    I_filtered_10b[473] = 10'h3A6;
    I_filtered_10b[472] = 10'h3C8;
    I_filtered_10b[471] = 10'h3EF;
    I_filtered_10b[470] = 10'h00F;
    I_filtered_10b[469] = 10'h032;
    I_filtered_10b[468] = 10'h050;
    I_filtered_10b[467] = 10'h06A;
    I_filtered_10b[466] = 10'h07F;
    I_filtered_10b[465] = 10'h090;
    I_filtered_10b[464] = 10'h099;
    I_filtered_10b[463] = 10'h09F;
    I_filtered_10b[462] = 10'h0A5;
    I_filtered_10b[461] = 10'h0A5;
    I_filtered_10b[460] = 10'h0A4;
    I_filtered_10b[459] = 10'h0A5;
    I_filtered_10b[458] = 10'h0A6;
    I_filtered_10b[457] = 10'h0A6;
    I_filtered_10b[456] = 10'h0AB;
    I_filtered_10b[455] = 10'h0AE;
    I_filtered_10b[454] = 10'h0B4;
    I_filtered_10b[453] = 10'h0B8;
    I_filtered_10b[452] = 10'h0BC;
    I_filtered_10b[451] = 10'h0C0;
    I_filtered_10b[450] = 10'h0C2;
    I_filtered_10b[449] = 10'h0C2;
    I_filtered_10b[448] = 10'h0BE;
    I_filtered_10b[447] = 10'h0BA;
    I_filtered_10b[446] = 10'h0B3;
    I_filtered_10b[445] = 10'h0AE;
    I_filtered_10b[444] = 10'h0A7;
    I_filtered_10b[443] = 10'h09E;
    I_filtered_10b[442] = 10'h099;
    I_filtered_10b[441] = 10'h092;
    I_filtered_10b[440] = 10'h08E;
    I_filtered_10b[439] = 10'h086;
    I_filtered_10b[438] = 10'h081;
    I_filtered_10b[437] = 10'h07B;
    I_filtered_10b[436] = 10'h076;
    I_filtered_10b[435] = 10'h074;
    I_filtered_10b[434] = 10'h070;
    I_filtered_10b[433] = 10'h06F;
    I_filtered_10b[432] = 10'h06B;
    I_filtered_10b[431] = 10'h06C;
    I_filtered_10b[430] = 10'h06C;
    I_filtered_10b[429] = 10'h06A;
    I_filtered_10b[428] = 10'h06B;
    I_filtered_10b[427] = 10'h06A;
    I_filtered_10b[426] = 10'h065;
    I_filtered_10b[425] = 10'h05F;
    I_filtered_10b[424] = 10'h059;
    I_filtered_10b[423] = 10'h04C;
    I_filtered_10b[422] = 10'h03B;
    I_filtered_10b[421] = 10'h026;
    I_filtered_10b[420] = 10'h00D;
    I_filtered_10b[419] = 10'h3EF;
    I_filtered_10b[418] = 10'h3D0;
    I_filtered_10b[417] = 10'h3AE;
    I_filtered_10b[416] = 10'h38D;
    I_filtered_10b[415] = 10'h372;
    I_filtered_10b[414] = 10'h35C;
    I_filtered_10b[413] = 10'h34F;
    I_filtered_10b[412] = 10'h349;
    I_filtered_10b[411] = 10'h34F;
    I_filtered_10b[410] = 10'h35F;
    I_filtered_10b[409] = 10'h378;
    I_filtered_10b[408] = 10'h397;
    I_filtered_10b[407] = 10'h3BE;
    I_filtered_10b[406] = 10'h3EA;
    I_filtered_10b[405] = 10'h014;
    I_filtered_10b[404] = 10'h03D;
    I_filtered_10b[403] = 10'h061;
    I_filtered_10b[402] = 10'h07C;
    I_filtered_10b[401] = 10'h092;
    I_filtered_10b[400] = 10'h0A0;
    I_filtered_10b[399] = 10'h0A5;
    I_filtered_10b[398] = 10'h0A2;
    I_filtered_10b[397] = 10'h09E;
    I_filtered_10b[396] = 10'h096;
    I_filtered_10b[395] = 10'h089;
    I_filtered_10b[394] = 10'h07F;
    I_filtered_10b[393] = 10'h073;
    I_filtered_10b[392] = 10'h06C;
    I_filtered_10b[391] = 10'h068;
    I_filtered_10b[390] = 10'h064;
    I_filtered_10b[389] = 10'h064;
    I_filtered_10b[388] = 10'h063;
    I_filtered_10b[387] = 10'h060;
    I_filtered_10b[386] = 10'h05F;
    I_filtered_10b[385] = 10'h05A;
    I_filtered_10b[384] = 10'h04F;
    I_filtered_10b[383] = 10'h03E;
    I_filtered_10b[382] = 10'h02C;
    I_filtered_10b[381] = 10'h011;
    I_filtered_10b[380] = 10'h3F6;
    I_filtered_10b[379] = 10'h3DA;
    I_filtered_10b[378] = 10'h3B8;
    I_filtered_10b[377] = 10'h39D;
    I_filtered_10b[376] = 10'h382;
    I_filtered_10b[375] = 10'h36E;
    I_filtered_10b[374] = 10'h35E;
    I_filtered_10b[373] = 10'h355;
    I_filtered_10b[372] = 10'h353;
    I_filtered_10b[371] = 10'h359;
    I_filtered_10b[370] = 10'h36A;
    I_filtered_10b[369] = 10'h37E;
    I_filtered_10b[368] = 10'h399;
    I_filtered_10b[367] = 10'h3B5;
    I_filtered_10b[366] = 10'h3D5;
    I_filtered_10b[365] = 10'h3F4;
    I_filtered_10b[364] = 10'h00E;
    I_filtered_10b[363] = 10'h025;
    I_filtered_10b[362] = 10'h037;
    I_filtered_10b[361] = 10'h041;
    I_filtered_10b[360] = 10'h044;
    I_filtered_10b[359] = 10'h041;
    I_filtered_10b[358] = 10'h034;
    I_filtered_10b[357] = 10'h01F;
    I_filtered_10b[356] = 10'h004;
    I_filtered_10b[355] = 10'h3E4;
    I_filtered_10b[354] = 10'h3C0;
    I_filtered_10b[353] = 10'h39A;
    I_filtered_10b[352] = 10'h374;
    I_filtered_10b[351] = 10'h353;
    I_filtered_10b[350] = 10'h334;
    I_filtered_10b[349] = 10'h31E;
    I_filtered_10b[348] = 10'h312;
    I_filtered_10b[347] = 10'h310;
    I_filtered_10b[346] = 10'h316;
    I_filtered_10b[345] = 10'h329;
    I_filtered_10b[344] = 10'h346;
    I_filtered_10b[343] = 10'h36D;
    I_filtered_10b[342] = 10'h399;
    I_filtered_10b[341] = 10'h3CE;
    I_filtered_10b[340] = 10'h002;
    I_filtered_10b[339] = 10'h036;
    I_filtered_10b[338] = 10'h067;
    I_filtered_10b[337] = 10'h08D;
    I_filtered_10b[336] = 10'h0AC;
    I_filtered_10b[335] = 10'h0BE;
    I_filtered_10b[334] = 10'h0C3;
    I_filtered_10b[333] = 10'h0BB;
    I_filtered_10b[332] = 10'h0AA;
    I_filtered_10b[331] = 10'h08E;
    I_filtered_10b[330] = 10'h06B;
    I_filtered_10b[329] = 10'h043;
    I_filtered_10b[328] = 10'h017;
    I_filtered_10b[327] = 10'h3EF;
    I_filtered_10b[326] = 10'h3C8;
    I_filtered_10b[325] = 10'h3A7;
    I_filtered_10b[324] = 10'h38C;
    I_filtered_10b[323] = 10'h376;
    I_filtered_10b[322] = 10'h367;
    I_filtered_10b[321] = 10'h361;
    I_filtered_10b[320] = 10'h35E;
    I_filtered_10b[319] = 10'h35D;
    I_filtered_10b[318] = 10'h361;
    I_filtered_10b[317] = 10'h369;
    I_filtered_10b[316] = 10'h36E;
    I_filtered_10b[315] = 10'h373;
    I_filtered_10b[314] = 10'h378;
    I_filtered_10b[313] = 10'h37A;
    I_filtered_10b[312] = 10'h37D;
    I_filtered_10b[311] = 10'h37F;
    I_filtered_10b[310] = 10'h380;
    I_filtered_10b[309] = 10'h381;
    I_filtered_10b[308] = 10'h37F;
    I_filtered_10b[307] = 10'h380;
    I_filtered_10b[306] = 10'h37E;
    I_filtered_10b[305] = 10'h37D;
    I_filtered_10b[304] = 10'h37A;
    I_filtered_10b[303] = 10'h378;
    I_filtered_10b[302] = 10'h376;
    I_filtered_10b[301] = 10'h372;
    I_filtered_10b[300] = 10'h36E;
    I_filtered_10b[299] = 10'h36A;
    I_filtered_10b[298] = 10'h365;
    I_filtered_10b[297] = 10'h362;
    I_filtered_10b[296] = 10'h364;
    I_filtered_10b[295] = 10'h367;
    I_filtered_10b[294] = 10'h36D;
    I_filtered_10b[293] = 10'h37A;
    I_filtered_10b[292] = 10'h38B;
    I_filtered_10b[291] = 10'h3A1;
    I_filtered_10b[290] = 10'h3BA;
    I_filtered_10b[289] = 10'h3D7;
    I_filtered_10b[288] = 10'h3F2;
    I_filtered_10b[287] = 10'h012;
    I_filtered_10b[286] = 10'h02E;
    I_filtered_10b[285] = 10'h04A;
    I_filtered_10b[284] = 10'h05E;
    I_filtered_10b[283] = 10'h06E;
    I_filtered_10b[282] = 10'h077;
    I_filtered_10b[281] = 10'h079;
    I_filtered_10b[280] = 10'h073;
    I_filtered_10b[279] = 10'h062;
    I_filtered_10b[278] = 10'h04D;
    I_filtered_10b[277] = 10'h031;
    I_filtered_10b[276] = 10'h013;
    I_filtered_10b[275] = 10'h3F1;
    I_filtered_10b[274] = 10'h3D1;
    I_filtered_10b[273] = 10'h3B5;
    I_filtered_10b[272] = 10'h39D;
    I_filtered_10b[271] = 10'h38B;
    I_filtered_10b[270] = 10'h383;
    I_filtered_10b[269] = 10'h383;
    I_filtered_10b[268] = 10'h38A;
    I_filtered_10b[267] = 10'h39B;
    I_filtered_10b[266] = 10'h3B4;
    I_filtered_10b[265] = 10'h3D5;
    I_filtered_10b[264] = 10'h3FA;
    I_filtered_10b[263] = 10'h023;
    I_filtered_10b[262] = 10'h04B;
    I_filtered_10b[261] = 10'h075;
    I_filtered_10b[260] = 10'h099;
    I_filtered_10b[259] = 10'h0BB;
    I_filtered_10b[258] = 10'h0D4;
    I_filtered_10b[257] = 10'h0E4;
    I_filtered_10b[256] = 10'h0EA;
    I_filtered_10b[255] = 10'h0E9;
    I_filtered_10b[254] = 10'h0DE;
    I_filtered_10b[253] = 10'h0C9;
    I_filtered_10b[252] = 10'h0AC;
    I_filtered_10b[251] = 10'h08B;
    I_filtered_10b[250] = 10'h066;
    I_filtered_10b[249] = 10'h040;
    I_filtered_10b[248] = 10'h01B;
    I_filtered_10b[247] = 10'h3FA;
    I_filtered_10b[246] = 10'h3DD;
    I_filtered_10b[245] = 10'h3C7;
    I_filtered_10b[244] = 10'h3BA;
    I_filtered_10b[243] = 10'h3B6;
    I_filtered_10b[242] = 10'h3BA;
    I_filtered_10b[241] = 10'h3C7;
    I_filtered_10b[240] = 10'h3DD;
    I_filtered_10b[239] = 10'h3FA;
    I_filtered_10b[238] = 10'h01B;
    I_filtered_10b[237] = 10'h041;
    I_filtered_10b[236] = 10'h068;
    I_filtered_10b[235] = 10'h08D;
    I_filtered_10b[234] = 10'h0AF;
    I_filtered_10b[233] = 10'h0CB;
    I_filtered_10b[232] = 10'h0E0;
    I_filtered_10b[231] = 10'h0EA;
    I_filtered_10b[230] = 10'h0EA;
    I_filtered_10b[229] = 10'h0E2;
    I_filtered_10b[228] = 10'h0D1;
    I_filtered_10b[227] = 10'h0B8;
    I_filtered_10b[226] = 10'h096;
    I_filtered_10b[225] = 10'h073;
    I_filtered_10b[224] = 10'h04A;
    I_filtered_10b[223] = 10'h025;
    I_filtered_10b[222] = 10'h3FF;
    I_filtered_10b[221] = 10'h3DD;
    I_filtered_10b[220] = 10'h3BF;
    I_filtered_10b[219] = 10'h3A8;
    I_filtered_10b[218] = 10'h397;
    I_filtered_10b[217] = 10'h38F;
    I_filtered_10b[216] = 10'h38C;
    I_filtered_10b[215] = 10'h38D;
    I_filtered_10b[214] = 10'h396;
    I_filtered_10b[213] = 10'h3A3;
    I_filtered_10b[212] = 10'h3B1;
    I_filtered_10b[211] = 10'h3BF;
    I_filtered_10b[210] = 10'h3CF;
    I_filtered_10b[209] = 10'h3DC;
    I_filtered_10b[208] = 10'h3E8;
    I_filtered_10b[207] = 10'h3F1;
    I_filtered_10b[206] = 10'h3F8;
    I_filtered_10b[205] = 10'h3FB;
    I_filtered_10b[204] = 10'h3F8;
    I_filtered_10b[203] = 10'h3F6;
    I_filtered_10b[202] = 10'h3ED;
    I_filtered_10b[201] = 10'h3E3;
    I_filtered_10b[200] = 10'h3D5;
    I_filtered_10b[199] = 10'h3C6;
    I_filtered_10b[198] = 10'h3B5;
    I_filtered_10b[197] = 10'h3A4;
    I_filtered_10b[196] = 10'h391;
    I_filtered_10b[195] = 10'h381;
    I_filtered_10b[194] = 10'h36F;
    I_filtered_10b[193] = 10'h363;
    I_filtered_10b[192] = 10'h35D;
    I_filtered_10b[191] = 10'h35B;
    I_filtered_10b[190] = 10'h35E;
    I_filtered_10b[189] = 10'h369;
    I_filtered_10b[188] = 10'h37C;
    I_filtered_10b[187] = 10'h395;
    I_filtered_10b[186] = 10'h3B2;
    I_filtered_10b[185] = 10'h3D6;
    I_filtered_10b[184] = 10'h3FC;
    I_filtered_10b[183] = 10'h020;
    I_filtered_10b[182] = 10'h044;
    I_filtered_10b[181] = 10'h05F;
    I_filtered_10b[180] = 10'h075;
    I_filtered_10b[179] = 10'h081;
    I_filtered_10b[178] = 10'h083;
    I_filtered_10b[177] = 10'h07A;
    I_filtered_10b[176] = 10'h068;
    I_filtered_10b[175] = 10'h04E;
    I_filtered_10b[174] = 10'h02E;
    I_filtered_10b[173] = 10'h008;
    I_filtered_10b[172] = 10'h3DF;
    I_filtered_10b[171] = 10'h3BA;
    I_filtered_10b[170] = 10'h394;
    I_filtered_10b[169] = 10'h375;
    I_filtered_10b[168] = 10'h35A;
    I_filtered_10b[167] = 10'h345;
    I_filtered_10b[166] = 10'h335;
    I_filtered_10b[165] = 10'h32E;
    I_filtered_10b[164] = 10'h329;
    I_filtered_10b[163] = 10'h327;
    I_filtered_10b[162] = 10'h32A;
    I_filtered_10b[161] = 10'h331;
    I_filtered_10b[160] = 10'h336;
    I_filtered_10b[159] = 10'h33A;
    I_filtered_10b[158] = 10'h33E;
    I_filtered_10b[157] = 10'h341;
    I_filtered_10b[156] = 10'h344;
    I_filtered_10b[155] = 10'h347;
    I_filtered_10b[154] = 10'h349;
    I_filtered_10b[153] = 10'h34C;
    I_filtered_10b[152] = 10'h34C;
    I_filtered_10b[151] = 10'h34F;
    I_filtered_10b[150] = 10'h34E;
    I_filtered_10b[149] = 10'h34C;
    I_filtered_10b[148] = 10'h34A;
    I_filtered_10b[147] = 10'h345;
    I_filtered_10b[146] = 10'h33F;
    I_filtered_10b[145] = 10'h334;
    I_filtered_10b[144] = 10'h32C;
    I_filtered_10b[143] = 10'h322;
    I_filtered_10b[142] = 10'h31A;
    I_filtered_10b[141] = 10'h315;
    I_filtered_10b[140] = 10'h31A;
    I_filtered_10b[139] = 10'h322;
    I_filtered_10b[138] = 10'h331;
    I_filtered_10b[137] = 10'h34A;
    I_filtered_10b[136] = 10'h368;
    I_filtered_10b[135] = 10'h38F;
    I_filtered_10b[134] = 10'h3B9;
    I_filtered_10b[133] = 10'h3EB;
    I_filtered_10b[132] = 10'h016;
    I_filtered_10b[131] = 10'h048;
    I_filtered_10b[130] = 10'h074;
    I_filtered_10b[129] = 10'h09C;
    I_filtered_10b[128] = 10'h0BB;
    I_filtered_10b[127] = 10'h0D5;
    I_filtered_10b[126] = 10'h0E4;
    I_filtered_10b[125] = 10'h0EB;
    I_filtered_10b[124] = 10'h0ED;
    I_filtered_10b[123] = 10'h0E3;
    I_filtered_10b[122] = 10'h0D7;
    I_filtered_10b[121] = 10'h0C5;
    I_filtered_10b[120] = 10'h0B6;
    I_filtered_10b[119] = 10'h0A3;
    I_filtered_10b[118] = 10'h093;
    I_filtered_10b[117] = 10'h088;
    I_filtered_10b[116] = 10'h07E;
    I_filtered_10b[115] = 10'h078;
    I_filtered_10b[114] = 10'h073;
    I_filtered_10b[113] = 10'h075;
    I_filtered_10b[112] = 10'h075;
    I_filtered_10b[111] = 10'h07A;
    I_filtered_10b[110] = 10'h081;
    I_filtered_10b[109] = 10'h08B;
    I_filtered_10b[108] = 10'h095;
    I_filtered_10b[107] = 10'h0A2;
    I_filtered_10b[106] = 10'h0B0;
    I_filtered_10b[105] = 10'h0BE;
    I_filtered_10b[104] = 10'h0CB;
    I_filtered_10b[103] = 10'h0D9;
    I_filtered_10b[102] = 10'h0E2;
    I_filtered_10b[101] = 10'h0E2;
    I_filtered_10b[100] = 10'h0DE;
    I_filtered_10b[99] = 10'h0D5;
    I_filtered_10b[98] = 10'h0C1;
    I_filtered_10b[97] = 10'h0A7;
    I_filtered_10b[96] = 10'h084;
    I_filtered_10b[95] = 10'h05D;
    I_filtered_10b[94] = 10'h02E;
    I_filtered_10b[93] = 10'h001;
    I_filtered_10b[92] = 10'h3D1;
    I_filtered_10b[91] = 10'h3A5;
    I_filtered_10b[90] = 10'h37F;
    I_filtered_10b[89] = 10'h361;
    I_filtered_10b[88] = 10'h34D;
    I_filtered_10b[87] = 10'h343;
    I_filtered_10b[86] = 10'h346;
    I_filtered_10b[85] = 10'h351;
    I_filtered_10b[84] = 10'h368;
    I_filtered_10b[83] = 10'h385;
    I_filtered_10b[82] = 10'h3A8;
    I_filtered_10b[81] = 10'h3CE;
    I_filtered_10b[80] = 10'h3F4;
    I_filtered_10b[79] = 10'h016;
    I_filtered_10b[78] = 10'h034;
    I_filtered_10b[77] = 10'h04B;
    I_filtered_10b[76] = 10'h05D;
    I_filtered_10b[75] = 10'h069;
    I_filtered_10b[74] = 10'h06B;
    I_filtered_10b[73] = 10'h06A;
    I_filtered_10b[72] = 10'h066;
    I_filtered_10b[71] = 10'h05E;
    I_filtered_10b[70] = 10'h052;
    I_filtered_10b[69] = 10'h048;
    I_filtered_10b[68] = 10'h03C;
    I_filtered_10b[67] = 10'h033;
    I_filtered_10b[66] = 10'h02B;
    I_filtered_10b[65] = 10'h023;
    I_filtered_10b[64] = 10'h01C;
    I_filtered_10b[63] = 10'h018;
    I_filtered_10b[62] = 10'h014;
    I_filtered_10b[61] = 10'h014;
    I_filtered_10b[60] = 10'h012;
    I_filtered_10b[59] = 10'h012;
    I_filtered_10b[58] = 10'h013;
    I_filtered_10b[57] = 10'h016;
    I_filtered_10b[56] = 10'h018;
    I_filtered_10b[55] = 10'h01C;
    I_filtered_10b[54] = 10'h020;
    I_filtered_10b[53] = 10'h024;
    I_filtered_10b[52] = 10'h029;
    I_filtered_10b[51] = 10'h02D;
    I_filtered_10b[50] = 10'h030;
    I_filtered_10b[49] = 10'h02F;
    I_filtered_10b[48] = 10'h02C;
    I_filtered_10b[47] = 10'h026;
    I_filtered_10b[46] = 10'h01B;
    I_filtered_10b[45] = 10'h00E;
    I_filtered_10b[44] = 10'h3FD;
    I_filtered_10b[43] = 10'h3EA;
    I_filtered_10b[42] = 10'h3D2;
    I_filtered_10b[41] = 10'h3BC;
    I_filtered_10b[40] = 10'h3A3;
    I_filtered_10b[39] = 10'h38D;
    I_filtered_10b[38] = 10'h37A;
    I_filtered_10b[37] = 10'h36C;
    I_filtered_10b[36] = 10'h362;
    I_filtered_10b[35] = 10'h35E;
    I_filtered_10b[34] = 10'h360;
    I_filtered_10b[33] = 10'h368;
    I_filtered_10b[32] = 10'h375;
    I_filtered_10b[31] = 10'h385;
    I_filtered_10b[30] = 10'h399;
    I_filtered_10b[29] = 10'h3AF;
    I_filtered_10b[28] = 10'h3C4;
    I_filtered_10b[27] = 10'h3D9;
    I_filtered_10b[26] = 10'h3EA;
    I_filtered_10b[25] = 10'h3F8;
    I_filtered_10b[24] = 10'h003;
    I_filtered_10b[23] = 10'h00C;
    I_filtered_10b[22] = 10'h00F;
    I_filtered_10b[21] = 10'h010;
    I_filtered_10b[20] = 10'h010;
    I_filtered_10b[19] = 10'h00D;
    I_filtered_10b[18] = 10'h009;
    I_filtered_10b[17] = 10'h006;
    I_filtered_10b[16] = 10'h002;
    I_filtered_10b[15] = 10'h3FF;
    I_filtered_10b[14] = 10'h3FE;
    I_filtered_10b[13] = 10'h3FC;
    I_filtered_10b[12] = 10'h3FC;
    I_filtered_10b[11] = 10'h3FC;
    I_filtered_10b[10] = 10'h3FE;
    I_filtered_10b[9] = 10'h000;
    I_filtered_10b[8] = 10'h001;
    I_filtered_10b[7] = 10'h002;
    I_filtered_10b[6] = 10'h002;
    I_filtered_10b[5] = 10'h004;
    I_filtered_10b[4] = 10'h002;
    I_filtered_10b[3] = 10'h002;
    I_filtered_10b[2] = 10'h001;
    I_filtered_10b[1] = 10'h000;
    I_filtered_10b[0] = 10'h000;


// Q Channel 10b Expected output
    Q_filtered_10b[1733] = 10'h000;
    Q_filtered_10b[1732] = 10'h000;
    Q_filtered_10b[1731] = 10'h000;
    Q_filtered_10b[1730] = 10'h000;
    Q_filtered_10b[1729] = 10'h000;
    Q_filtered_10b[1728] = 10'h000;
    Q_filtered_10b[1727] = 10'h000;
    Q_filtered_10b[1726] = 10'h000;
    Q_filtered_10b[1725] = 10'h000;
    Q_filtered_10b[1724] = 10'h000;
    Q_filtered_10b[1723] = 10'h000;
    Q_filtered_10b[1722] = 10'h000;
    Q_filtered_10b[1721] = 10'h000;
    Q_filtered_10b[1720] = 10'h000;
    Q_filtered_10b[1719] = 10'h001;
    Q_filtered_10b[1718] = 10'h002;
    Q_filtered_10b[1717] = 10'h002;
    Q_filtered_10b[1716] = 10'h004;
    Q_filtered_10b[1715] = 10'h002;
    Q_filtered_10b[1714] = 10'h002;
    Q_filtered_10b[1713] = 10'h001;
    Q_filtered_10b[1712] = 10'h000;
    Q_filtered_10b[1711] = 10'h3FE;
    Q_filtered_10b[1710] = 10'h3FC;
    Q_filtered_10b[1709] = 10'h3FC;
    Q_filtered_10b[1708] = 10'h3FC;
    Q_filtered_10b[1707] = 10'h3FE;
    Q_filtered_10b[1706] = 10'h3FE;
    Q_filtered_10b[1705] = 10'h001;
    Q_filtered_10b[1704] = 10'h005;
    Q_filtered_10b[1703] = 10'h006;
    Q_filtered_10b[1702] = 10'h00B;
    Q_filtered_10b[1701] = 10'h00D;
    Q_filtered_10b[1700] = 10'h00E;
    Q_filtered_10b[1699] = 10'h00E;
    Q_filtered_10b[1698] = 10'h00B;
    Q_filtered_10b[1697] = 10'h005;
    Q_filtered_10b[1696] = 10'h3FB;
    Q_filtered_10b[1695] = 10'h3EE;
    Q_filtered_10b[1694] = 10'h3DD;
    Q_filtered_10b[1693] = 10'h3CA;
    Q_filtered_10b[1692] = 10'h3B4;
    Q_filtered_10b[1691] = 10'h39F;
    Q_filtered_10b[1690] = 10'h38C;
    Q_filtered_10b[1689] = 10'h37C;
    Q_filtered_10b[1688] = 10'h36F;
    Q_filtered_10b[1687] = 10'h369;
    Q_filtered_10b[1686] = 10'h369;
    Q_filtered_10b[1685] = 10'h36F;
    Q_filtered_10b[1684] = 10'h37D;
    Q_filtered_10b[1683] = 10'h38E;
    Q_filtered_10b[1682] = 10'h3A4;
    Q_filtered_10b[1681] = 10'h3BD;
    Q_filtered_10b[1680] = 10'h3D8;
    Q_filtered_10b[1679] = 10'h3F1;
    Q_filtered_10b[1678] = 10'h00A;
    Q_filtered_10b[1677] = 10'h020;
    Q_filtered_10b[1676] = 10'h033;
    Q_filtered_10b[1675] = 10'h041;
    Q_filtered_10b[1674] = 10'h04E;
    Q_filtered_10b[1673] = 10'h055;
    Q_filtered_10b[1672] = 10'h05C;
    Q_filtered_10b[1671] = 10'h060;
    Q_filtered_10b[1670] = 10'h061;
    Q_filtered_10b[1669] = 10'h061;
    Q_filtered_10b[1668] = 10'h064;
    Q_filtered_10b[1667] = 10'h066;
    Q_filtered_10b[1666] = 10'h067;
    Q_filtered_10b[1665] = 10'h06B;
    Q_filtered_10b[1664] = 10'h06F;
    Q_filtered_10b[1663] = 10'h071;
    Q_filtered_10b[1662] = 10'h074;
    Q_filtered_10b[1661] = 10'h077;
    Q_filtered_10b[1660] = 10'h078;
    Q_filtered_10b[1659] = 10'h079;
    Q_filtered_10b[1658] = 10'h079;
    Q_filtered_10b[1657] = 10'h079;
    Q_filtered_10b[1656] = 10'h07A;
    Q_filtered_10b[1655] = 10'h07C;
    Q_filtered_10b[1654] = 10'h07D;
    Q_filtered_10b[1653] = 10'h081;
    Q_filtered_10b[1652] = 10'h086;
    Q_filtered_10b[1651] = 10'h088;
    Q_filtered_10b[1650] = 10'h08F;
    Q_filtered_10b[1649] = 10'h093;
    Q_filtered_10b[1648] = 10'h093;
    Q_filtered_10b[1647] = 10'h08E;
    Q_filtered_10b[1646] = 10'h089;
    Q_filtered_10b[1645] = 10'h07A;
    Q_filtered_10b[1644] = 10'h067;
    Q_filtered_10b[1643] = 10'h04F;
    Q_filtered_10b[1642] = 10'h031;
    Q_filtered_10b[1641] = 10'h011;
    Q_filtered_10b[1640] = 10'h3F0;
    Q_filtered_10b[1639] = 10'h3CB;
    Q_filtered_10b[1638] = 10'h3AC;
    Q_filtered_10b[1637] = 10'h38D;
    Q_filtered_10b[1636] = 10'h376;
    Q_filtered_10b[1635] = 10'h364;
    Q_filtered_10b[1634] = 10'h35C;
    Q_filtered_10b[1633] = 10'h359;
    Q_filtered_10b[1632] = 10'h362;
    Q_filtered_10b[1631] = 10'h376;
    Q_filtered_10b[1630] = 10'h38F;
    Q_filtered_10b[1629] = 10'h3AE;
    Q_filtered_10b[1628] = 10'h3D1;
    Q_filtered_10b[1627] = 10'h3F9;
    Q_filtered_10b[1626] = 10'h01D;
    Q_filtered_10b[1625] = 10'h03C;
    Q_filtered_10b[1624] = 10'h057;
    Q_filtered_10b[1623] = 10'h06B;
    Q_filtered_10b[1622] = 10'h076;
    Q_filtered_10b[1621] = 10'h076;
    Q_filtered_10b[1620] = 10'h071;
    Q_filtered_10b[1619] = 10'h061;
    Q_filtered_10b[1618] = 10'h04A;
    Q_filtered_10b[1617] = 10'h02A;
    Q_filtered_10b[1616] = 10'h008;
    Q_filtered_10b[1615] = 10'h3E0;
    Q_filtered_10b[1614] = 10'h3B7;
    Q_filtered_10b[1613] = 10'h392;
    Q_filtered_10b[1612] = 10'h36F;
    Q_filtered_10b[1611] = 10'h352;
    Q_filtered_10b[1610] = 10'h33C;
    Q_filtered_10b[1609] = 10'h32F;
    Q_filtered_10b[1608] = 10'h32E;
    Q_filtered_10b[1607] = 10'h331;
    Q_filtered_10b[1606] = 10'h33F;
    Q_filtered_10b[1605] = 10'h352;
    Q_filtered_10b[1604] = 10'h36D;
    Q_filtered_10b[1603] = 10'h387;
    Q_filtered_10b[1602] = 10'h3A8;
    Q_filtered_10b[1601] = 10'h3C8;
    Q_filtered_10b[1600] = 10'h3E3;
    Q_filtered_10b[1599] = 10'h3FF;
    Q_filtered_10b[1598] = 10'h011;
    Q_filtered_10b[1597] = 10'h021;
    Q_filtered_10b[1596] = 10'h02A;
    Q_filtered_10b[1595] = 10'h02D;
    Q_filtered_10b[1594] = 10'h02B;
    Q_filtered_10b[1593] = 10'h028;
    Q_filtered_10b[1592] = 10'h025;
    Q_filtered_10b[1591] = 10'h01E;
    Q_filtered_10b[1590] = 10'h01D;
    Q_filtered_10b[1589] = 10'h01A;
    Q_filtered_10b[1588] = 10'h01B;
    Q_filtered_10b[1587] = 10'h01F;
    Q_filtered_10b[1586] = 10'h021;
    Q_filtered_10b[1585] = 10'h027;
    Q_filtered_10b[1584] = 10'h02A;
    Q_filtered_10b[1583] = 10'h02C;
    Q_filtered_10b[1582] = 10'h02D;
    Q_filtered_10b[1581] = 10'h028;
    Q_filtered_10b[1580] = 10'h01E;
    Q_filtered_10b[1579] = 10'h00E;
    Q_filtered_10b[1578] = 10'h3FC;
    Q_filtered_10b[1577] = 10'h3E1;
    Q_filtered_10b[1576] = 10'h3C6;
    Q_filtered_10b[1575] = 10'h3A7;
    Q_filtered_10b[1574] = 10'h389;
    Q_filtered_10b[1573] = 10'h36F;
    Q_filtered_10b[1572] = 10'h359;
    Q_filtered_10b[1571] = 10'h348;
    Q_filtered_10b[1570] = 10'h33C;
    Q_filtered_10b[1569] = 10'h339;
    Q_filtered_10b[1568] = 10'h33A;
    Q_filtered_10b[1567] = 10'h343;
    Q_filtered_10b[1566] = 10'h351;
    Q_filtered_10b[1565] = 10'h364;
    Q_filtered_10b[1564] = 10'h378;
    Q_filtered_10b[1563] = 10'h390;
    Q_filtered_10b[1562] = 10'h3A7;
    Q_filtered_10b[1561] = 10'h3BC;
    Q_filtered_10b[1560] = 10'h3D0;
    Q_filtered_10b[1559] = 10'h3DD;
    Q_filtered_10b[1558] = 10'h3E8;
    Q_filtered_10b[1557] = 10'h3F0;
    Q_filtered_10b[1556] = 10'h3F4;
    Q_filtered_10b[1555] = 10'h3F5;
    Q_filtered_10b[1554] = 10'h3F7;
    Q_filtered_10b[1553] = 10'h3F8;
    Q_filtered_10b[1552] = 10'h3F8;
    Q_filtered_10b[1551] = 10'h3FC;
    Q_filtered_10b[1550] = 10'h3FD;
    Q_filtered_10b[1549] = 10'h001;
    Q_filtered_10b[1548] = 10'h009;
    Q_filtered_10b[1547] = 10'h00E;
    Q_filtered_10b[1546] = 10'h017;
    Q_filtered_10b[1545] = 10'h01C;
    Q_filtered_10b[1544] = 10'h022;
    Q_filtered_10b[1543] = 10'h027;
    Q_filtered_10b[1542] = 10'h029;
    Q_filtered_10b[1541] = 10'h026;
    Q_filtered_10b[1540] = 10'h01E;
    Q_filtered_10b[1539] = 10'h014;
    Q_filtered_10b[1538] = 10'h004;
    Q_filtered_10b[1537] = 10'h3F4;
    Q_filtered_10b[1536] = 10'h3DF;
    Q_filtered_10b[1535] = 10'h3CA;
    Q_filtered_10b[1534] = 10'h3BB;
    Q_filtered_10b[1533] = 10'h3AB;
    Q_filtered_10b[1532] = 10'h3A0;
    Q_filtered_10b[1531] = 10'h39A;
    Q_filtered_10b[1530] = 10'h39A;
    Q_filtered_10b[1529] = 10'h39E;
    Q_filtered_10b[1528] = 10'h3AA;
    Q_filtered_10b[1527] = 10'h3BB;
    Q_filtered_10b[1526] = 10'h3D2;
    Q_filtered_10b[1525] = 10'h3EC;
    Q_filtered_10b[1524] = 10'h009;
    Q_filtered_10b[1523] = 10'h027;
    Q_filtered_10b[1522] = 10'h045;
    Q_filtered_10b[1521] = 10'h05E;
    Q_filtered_10b[1520] = 10'h077;
    Q_filtered_10b[1519] = 10'h088;
    Q_filtered_10b[1518] = 10'h095;
    Q_filtered_10b[1517] = 10'h099;
    Q_filtered_10b[1516] = 10'h09A;
    Q_filtered_10b[1515] = 10'h092;
    Q_filtered_10b[1514] = 10'h084;
    Q_filtered_10b[1513] = 10'h070;
    Q_filtered_10b[1512] = 10'h05A;
    Q_filtered_10b[1511] = 10'h03F;
    Q_filtered_10b[1510] = 10'h021;
    Q_filtered_10b[1509] = 10'h008;
    Q_filtered_10b[1508] = 10'h3F0;
    Q_filtered_10b[1507] = 10'h3DE;
    Q_filtered_10b[1506] = 10'h3CF;
    Q_filtered_10b[1505] = 10'h3C8;
    Q_filtered_10b[1504] = 10'h3C8;
    Q_filtered_10b[1503] = 10'h3CE;
    Q_filtered_10b[1502] = 10'h3D9;
    Q_filtered_10b[1501] = 10'h3E8;
    Q_filtered_10b[1500] = 10'h3FC;
    Q_filtered_10b[1499] = 10'h010;
    Q_filtered_10b[1498] = 10'h027;
    Q_filtered_10b[1497] = 10'h03D;
    Q_filtered_10b[1496] = 10'h050;
    Q_filtered_10b[1495] = 10'h062;
    Q_filtered_10b[1494] = 10'h070;
    Q_filtered_10b[1493] = 10'h07A;
    Q_filtered_10b[1492] = 10'h082;
    Q_filtered_10b[1491] = 10'h083;
    Q_filtered_10b[1490] = 10'h085;
    Q_filtered_10b[1489] = 10'h084;
    Q_filtered_10b[1488] = 10'h083;
    Q_filtered_10b[1487] = 10'h07E;
    Q_filtered_10b[1486] = 10'h07F;
    Q_filtered_10b[1485] = 10'h07D;
    Q_filtered_10b[1484] = 10'h07D;
    Q_filtered_10b[1483] = 10'h07E;
    Q_filtered_10b[1482] = 10'h07E;
    Q_filtered_10b[1481] = 10'h07F;
    Q_filtered_10b[1480] = 10'h080;
    Q_filtered_10b[1479] = 10'h080;
    Q_filtered_10b[1478] = 10'h07E;
    Q_filtered_10b[1477] = 10'h07C;
    Q_filtered_10b[1476] = 10'h076;
    Q_filtered_10b[1475] = 10'h06F;
    Q_filtered_10b[1474] = 10'h067;
    Q_filtered_10b[1473] = 10'h05C;
    Q_filtered_10b[1472] = 10'h051;
    Q_filtered_10b[1471] = 10'h046;
    Q_filtered_10b[1470] = 10'h03A;
    Q_filtered_10b[1469] = 10'h02E;
    Q_filtered_10b[1468] = 10'h026;
    Q_filtered_10b[1467] = 10'h01E;
    Q_filtered_10b[1466] = 10'h017;
    Q_filtered_10b[1465] = 10'h011;
    Q_filtered_10b[1464] = 10'h00E;
    Q_filtered_10b[1463] = 10'h00A;
    Q_filtered_10b[1462] = 10'h009;
    Q_filtered_10b[1461] = 10'h006;
    Q_filtered_10b[1460] = 10'h003;
    Q_filtered_10b[1459] = 10'h000;
    Q_filtered_10b[1458] = 10'h3FD;
    Q_filtered_10b[1457] = 10'h3F8;
    Q_filtered_10b[1456] = 10'h3F3;
    Q_filtered_10b[1455] = 10'h3EC;
    Q_filtered_10b[1454] = 10'h3E7;
    Q_filtered_10b[1453] = 10'h3E2;
    Q_filtered_10b[1452] = 10'h3DE;
    Q_filtered_10b[1451] = 10'h3DC;
    Q_filtered_10b[1450] = 10'h3DD;
    Q_filtered_10b[1449] = 10'h3E2;
    Q_filtered_10b[1448] = 10'h3E7;
    Q_filtered_10b[1447] = 10'h3F0;
    Q_filtered_10b[1446] = 10'h3F8;
    Q_filtered_10b[1445] = 10'h003;
    Q_filtered_10b[1444] = 10'h00E;
    Q_filtered_10b[1443] = 10'h015;
    Q_filtered_10b[1442] = 10'h01E;
    Q_filtered_10b[1441] = 10'h023;
    Q_filtered_10b[1440] = 10'h027;
    Q_filtered_10b[1439] = 10'h027;
    Q_filtered_10b[1438] = 10'h026;
    Q_filtered_10b[1437] = 10'h021;
    Q_filtered_10b[1436] = 10'h018;
    Q_filtered_10b[1435] = 10'h00D;
    Q_filtered_10b[1434] = 10'h3FF;
    Q_filtered_10b[1433] = 10'h3ED;
    Q_filtered_10b[1432] = 10'h3DA;
    Q_filtered_10b[1431] = 10'h3C9;
    Q_filtered_10b[1430] = 10'h3B8;
    Q_filtered_10b[1429] = 10'h3AC;
    Q_filtered_10b[1428] = 10'h3A2;
    Q_filtered_10b[1427] = 10'h39E;
    Q_filtered_10b[1426] = 10'h3A0;
    Q_filtered_10b[1425] = 10'h3A6;
    Q_filtered_10b[1424] = 10'h3B1;
    Q_filtered_10b[1423] = 10'h3BE;
    Q_filtered_10b[1422] = 10'h3D0;
    Q_filtered_10b[1421] = 10'h3E2;
    Q_filtered_10b[1420] = 10'h3F5;
    Q_filtered_10b[1419] = 10'h005;
    Q_filtered_10b[1418] = 10'h015;
    Q_filtered_10b[1417] = 10'h024;
    Q_filtered_10b[1416] = 10'h031;
    Q_filtered_10b[1415] = 10'h03A;
    Q_filtered_10b[1414] = 10'h044;
    Q_filtered_10b[1413] = 10'h04A;
    Q_filtered_10b[1412] = 10'h053;
    Q_filtered_10b[1411] = 10'h05A;
    Q_filtered_10b[1410] = 10'h060;
    Q_filtered_10b[1409] = 10'h066;
    Q_filtered_10b[1408] = 10'h070;
    Q_filtered_10b[1407] = 10'h07B;
    Q_filtered_10b[1406] = 10'h084;
    Q_filtered_10b[1405] = 10'h08E;
    Q_filtered_10b[1404] = 10'h098;
    Q_filtered_10b[1403] = 10'h09F;
    Q_filtered_10b[1402] = 10'h0A5;
    Q_filtered_10b[1401] = 10'h0AA;
    Q_filtered_10b[1400] = 10'h0AC;
    Q_filtered_10b[1399] = 10'h0AD;
    Q_filtered_10b[1398] = 10'h0AC;
    Q_filtered_10b[1397] = 10'h0AC;
    Q_filtered_10b[1396] = 10'h0AC;
    Q_filtered_10b[1395] = 10'h0AE;
    Q_filtered_10b[1394] = 10'h0B0;
    Q_filtered_10b[1393] = 10'h0B5;
    Q_filtered_10b[1392] = 10'h0BB;
    Q_filtered_10b[1391] = 10'h0BE;
    Q_filtered_10b[1390] = 10'h0C5;
    Q_filtered_10b[1389] = 10'h0C9;
    Q_filtered_10b[1388] = 10'h0C8;
    Q_filtered_10b[1387] = 10'h0C2;
    Q_filtered_10b[1386] = 10'h0B9;
    Q_filtered_10b[1385] = 10'h0A6;
    Q_filtered_10b[1384] = 10'h090;
    Q_filtered_10b[1383] = 10'h073;
    Q_filtered_10b[1382] = 10'h051;
    Q_filtered_10b[1381] = 10'h02C;
    Q_filtered_10b[1380] = 10'h008;
    Q_filtered_10b[1379] = 10'h3E0;
    Q_filtered_10b[1378] = 10'h3BD;
    Q_filtered_10b[1377] = 10'h39B;
    Q_filtered_10b[1376] = 10'h383;
    Q_filtered_10b[1375] = 10'h36D;
    Q_filtered_10b[1374] = 10'h361;
    Q_filtered_10b[1373] = 10'h35B;
    Q_filtered_10b[1372] = 10'h35D;
    Q_filtered_10b[1371] = 10'h36A;
    Q_filtered_10b[1370] = 10'h37A;
    Q_filtered_10b[1369] = 10'h38E;
    Q_filtered_10b[1368] = 10'h3A5;
    Q_filtered_10b[1367] = 10'h3C1;
    Q_filtered_10b[1366] = 10'h3D7;
    Q_filtered_10b[1365] = 10'h3EA;
    Q_filtered_10b[1364] = 10'h3F8;
    Q_filtered_10b[1363] = 10'h003;
    Q_filtered_10b[1362] = 10'h007;
    Q_filtered_10b[1361] = 10'h004;
    Q_filtered_10b[1360] = 10'h3FE;
    Q_filtered_10b[1359] = 10'h3F2;
    Q_filtered_10b[1358] = 10'h3E4;
    Q_filtered_10b[1357] = 10'h3D0;
    Q_filtered_10b[1356] = 10'h3BC;
    Q_filtered_10b[1355] = 10'h3A4;
    Q_filtered_10b[1354] = 10'h38D;
    Q_filtered_10b[1353] = 10'h379;
    Q_filtered_10b[1352] = 10'h365;
    Q_filtered_10b[1351] = 10'h355;
    Q_filtered_10b[1350] = 10'h349;
    Q_filtered_10b[1349] = 10'h342;
    Q_filtered_10b[1348] = 10'h344;
    Q_filtered_10b[1347] = 10'h346;
    Q_filtered_10b[1346] = 10'h34E;
    Q_filtered_10b[1345] = 10'h357;
    Q_filtered_10b[1344] = 10'h365;
    Q_filtered_10b[1343] = 10'h370;
    Q_filtered_10b[1342] = 10'h37D;
    Q_filtered_10b[1341] = 10'h387;
    Q_filtered_10b[1340] = 10'h391;
    Q_filtered_10b[1339] = 10'h39B;
    Q_filtered_10b[1338] = 10'h3A2;
    Q_filtered_10b[1337] = 10'h3A8;
    Q_filtered_10b[1336] = 10'h3AF;
    Q_filtered_10b[1335] = 10'h3B6;
    Q_filtered_10b[1334] = 10'h3BC;
    Q_filtered_10b[1333] = 10'h3C6;
    Q_filtered_10b[1332] = 10'h3CF;
    Q_filtered_10b[1331] = 10'h3DB;
    Q_filtered_10b[1330] = 10'h3EA;
    Q_filtered_10b[1329] = 10'h3F8;
    Q_filtered_10b[1328] = 10'h005;
    Q_filtered_10b[1327] = 10'h016;
    Q_filtered_10b[1326] = 10'h025;
    Q_filtered_10b[1325] = 10'h035;
    Q_filtered_10b[1324] = 10'h040;
    Q_filtered_10b[1323] = 10'h04C;
    Q_filtered_10b[1322] = 10'h055;
    Q_filtered_10b[1321] = 10'h05D;
    Q_filtered_10b[1320] = 10'h060;
    Q_filtered_10b[1319] = 10'h05E;
    Q_filtered_10b[1318] = 10'h05C;
    Q_filtered_10b[1317] = 10'h057;
    Q_filtered_10b[1316] = 10'h053;
    Q_filtered_10b[1315] = 10'h04A;
    Q_filtered_10b[1314] = 10'h043;
    Q_filtered_10b[1313] = 10'h03F;
    Q_filtered_10b[1312] = 10'h03B;
    Q_filtered_10b[1311] = 10'h038;
    Q_filtered_10b[1310] = 10'h038;
    Q_filtered_10b[1309] = 10'h03A;
    Q_filtered_10b[1308] = 10'h03E;
    Q_filtered_10b[1307] = 10'h044;
    Q_filtered_10b[1306] = 10'h04D;
    Q_filtered_10b[1305] = 10'h059;
    Q_filtered_10b[1304] = 10'h067;
    Q_filtered_10b[1303] = 10'h078;
    Q_filtered_10b[1302] = 10'h08B;
    Q_filtered_10b[1301] = 10'h09C;
    Q_filtered_10b[1300] = 10'h0AC;
    Q_filtered_10b[1299] = 10'h0B8;
    Q_filtered_10b[1298] = 10'h0C2;
    Q_filtered_10b[1297] = 10'h0C6;
    Q_filtered_10b[1296] = 10'h0C2;
    Q_filtered_10b[1295] = 10'h0BA;
    Q_filtered_10b[1294] = 10'h0AC;
    Q_filtered_10b[1293] = 10'h09C;
    Q_filtered_10b[1292] = 10'h086;
    Q_filtered_10b[1291] = 10'h070;
    Q_filtered_10b[1290] = 10'h055;
    Q_filtered_10b[1289] = 10'h03E;
    Q_filtered_10b[1288] = 10'h028;
    Q_filtered_10b[1287] = 10'h011;
    Q_filtered_10b[1286] = 10'h003;
    Q_filtered_10b[1285] = 10'h3F7;
    Q_filtered_10b[1284] = 10'h3EB;
    Q_filtered_10b[1283] = 10'h3E4;
    Q_filtered_10b[1282] = 10'h3DF;
    Q_filtered_10b[1281] = 10'h3D6;
    Q_filtered_10b[1280] = 10'h3CE;
    Q_filtered_10b[1279] = 10'h3C4;
    Q_filtered_10b[1278] = 10'h3B3;
    Q_filtered_10b[1277] = 10'h3A4;
    Q_filtered_10b[1276] = 10'h391;
    Q_filtered_10b[1275] = 10'h379;
    Q_filtered_10b[1274] = 10'h366;
    Q_filtered_10b[1273] = 10'h34E;
    Q_filtered_10b[1272] = 10'h33E;
    Q_filtered_10b[1271] = 10'h332;
    Q_filtered_10b[1270] = 10'h32E;
    Q_filtered_10b[1269] = 10'h32F;
    Q_filtered_10b[1268] = 10'h33E;
    Q_filtered_10b[1267] = 10'h357;
    Q_filtered_10b[1266] = 10'h376;
    Q_filtered_10b[1265] = 10'h3A0;
    Q_filtered_10b[1264] = 10'h3CA;
    Q_filtered_10b[1263] = 10'h3FA;
    Q_filtered_10b[1262] = 10'h02B;
    Q_filtered_10b[1261] = 10'h052;
    Q_filtered_10b[1260] = 10'h078;
    Q_filtered_10b[1259] = 10'h094;
    Q_filtered_10b[1258] = 10'h0A8;
    Q_filtered_10b[1257] = 10'h0AF;
    Q_filtered_10b[1256] = 10'h0B0;
    Q_filtered_10b[1255] = 10'h0A3;
    Q_filtered_10b[1254] = 10'h08A;
    Q_filtered_10b[1253] = 10'h06A;
    Q_filtered_10b[1252] = 10'h044;
    Q_filtered_10b[1251] = 10'h01A;
    Q_filtered_10b[1250] = 10'h3EB;
    Q_filtered_10b[1249] = 10'h3BF;
    Q_filtered_10b[1248] = 10'h39B;
    Q_filtered_10b[1247] = 10'h379;
    Q_filtered_10b[1246] = 10'h360;
    Q_filtered_10b[1245] = 10'h352;
    Q_filtered_10b[1244] = 10'h351;
    Q_filtered_10b[1243] = 10'h355;
    Q_filtered_10b[1242] = 10'h368;
    Q_filtered_10b[1241] = 10'h383;
    Q_filtered_10b[1240] = 10'h3A9;
    Q_filtered_10b[1239] = 10'h3D2;
    Q_filtered_10b[1238] = 10'h004;
    Q_filtered_10b[1237] = 10'h039;
    Q_filtered_10b[1236] = 10'h068;
    Q_filtered_10b[1235] = 10'h094;
    Q_filtered_10b[1234] = 10'h0B8;
    Q_filtered_10b[1233] = 10'h0D4;
    Q_filtered_10b[1232] = 10'h0E3;
    Q_filtered_10b[1231] = 10'h0E3;
    Q_filtered_10b[1230] = 10'h0DA;
    Q_filtered_10b[1229] = 10'h0C5;
    Q_filtered_10b[1228] = 10'h0A9;
    Q_filtered_10b[1227] = 10'h082;
    Q_filtered_10b[1226] = 10'h05C;
    Q_filtered_10b[1225] = 10'h02F;
    Q_filtered_10b[1224] = 10'h005;
    Q_filtered_10b[1223] = 10'h3DF;
    Q_filtered_10b[1222] = 10'h3BB;
    Q_filtered_10b[1221] = 10'h39F;
    Q_filtered_10b[1220] = 10'h38A;
    Q_filtered_10b[1219] = 10'h378;
    Q_filtered_10b[1218] = 10'h372;
    Q_filtered_10b[1217] = 10'h36C;
    Q_filtered_10b[1216] = 10'h369;
    Q_filtered_10b[1215] = 10'h36A;
    Q_filtered_10b[1214] = 10'h36E;
    Q_filtered_10b[1213] = 10'h36A;
    Q_filtered_10b[1212] = 10'h36A;
    Q_filtered_10b[1211] = 10'h368;
    Q_filtered_10b[1210] = 10'h362;
    Q_filtered_10b[1209] = 10'h35E;
    Q_filtered_10b[1208] = 10'h358;
    Q_filtered_10b[1207] = 10'h354;
    Q_filtered_10b[1206] = 10'h350;
    Q_filtered_10b[1205] = 10'h34F;
    Q_filtered_10b[1204] = 10'h34F;
    Q_filtered_10b[1203] = 10'h354;
    Q_filtered_10b[1202] = 10'h35B;
    Q_filtered_10b[1201] = 10'h363;
    Q_filtered_10b[1200] = 10'h36F;
    Q_filtered_10b[1199] = 10'h37A;
    Q_filtered_10b[1198] = 10'h385;
    Q_filtered_10b[1197] = 10'h391;
    Q_filtered_10b[1196] = 10'h39B;
    Q_filtered_10b[1195] = 10'h3A1;
    Q_filtered_10b[1194] = 10'h3A7;
    Q_filtered_10b[1193] = 10'h3AE;
    Q_filtered_10b[1192] = 10'h3B6;
    Q_filtered_10b[1191] = 10'h3BB;
    Q_filtered_10b[1190] = 10'h3C5;
    Q_filtered_10b[1189] = 10'h3CE;
    Q_filtered_10b[1188] = 10'h3DB;
    Q_filtered_10b[1187] = 10'h3EA;
    Q_filtered_10b[1186] = 10'h3FB;
    Q_filtered_10b[1185] = 10'h00D;
    Q_filtered_10b[1184] = 10'h020;
    Q_filtered_10b[1183] = 10'h033;
    Q_filtered_10b[1182] = 10'h044;
    Q_filtered_10b[1181] = 10'h051;
    Q_filtered_10b[1180] = 10'h05B;
    Q_filtered_10b[1179] = 10'h060;
    Q_filtered_10b[1178] = 10'h060;
    Q_filtered_10b[1177] = 10'h05B;
    Q_filtered_10b[1176] = 10'h051;
    Q_filtered_10b[1175] = 10'h045;
    Q_filtered_10b[1174] = 10'h035;
    Q_filtered_10b[1173] = 10'h024;
    Q_filtered_10b[1172] = 10'h012;
    Q_filtered_10b[1171] = 10'h003;
    Q_filtered_10b[1170] = 10'h3F6;
    Q_filtered_10b[1169] = 10'h3EF;
    Q_filtered_10b[1168] = 10'h3E8;
    Q_filtered_10b[1167] = 10'h3E4;
    Q_filtered_10b[1166] = 10'h3E4;
    Q_filtered_10b[1165] = 10'h3E4;
    Q_filtered_10b[1164] = 10'h3E3;
    Q_filtered_10b[1163] = 10'h3E1;
    Q_filtered_10b[1162] = 10'h3DF;
    Q_filtered_10b[1161] = 10'h3D8;
    Q_filtered_10b[1160] = 10'h3D2;
    Q_filtered_10b[1159] = 10'h3C7;
    Q_filtered_10b[1158] = 10'h3BC;
    Q_filtered_10b[1157] = 10'h3B3;
    Q_filtered_10b[1156] = 10'h3A9;
    Q_filtered_10b[1155] = 10'h3A2;
    Q_filtered_10b[1154] = 10'h39F;
    Q_filtered_10b[1153] = 10'h3A0;
    Q_filtered_10b[1152] = 10'h3A5;
    Q_filtered_10b[1151] = 10'h3B1;
    Q_filtered_10b[1150] = 10'h3C1;
    Q_filtered_10b[1149] = 10'h3D5;
    Q_filtered_10b[1148] = 10'h3EF;
    Q_filtered_10b[1147] = 10'h00B;
    Q_filtered_10b[1146] = 10'h028;
    Q_filtered_10b[1145] = 10'h044;
    Q_filtered_10b[1144] = 10'h05D;
    Q_filtered_10b[1143] = 10'h070;
    Q_filtered_10b[1142] = 10'h080;
    Q_filtered_10b[1141] = 10'h08B;
    Q_filtered_10b[1140] = 10'h08E;
    Q_filtered_10b[1139] = 10'h08E;
    Q_filtered_10b[1138] = 10'h08A;
    Q_filtered_10b[1137] = 10'h083;
    Q_filtered_10b[1136] = 10'h07A;
    Q_filtered_10b[1135] = 10'h073;
    Q_filtered_10b[1134] = 10'h068;
    Q_filtered_10b[1133] = 10'h060;
    Q_filtered_10b[1132] = 10'h05C;
    Q_filtered_10b[1131] = 10'h056;
    Q_filtered_10b[1130] = 10'h058;
    Q_filtered_10b[1129] = 10'h057;
    Q_filtered_10b[1128] = 10'h056;
    Q_filtered_10b[1127] = 10'h055;
    Q_filtered_10b[1126] = 10'h054;
    Q_filtered_10b[1125] = 10'h04A;
    Q_filtered_10b[1124] = 10'h03C;
    Q_filtered_10b[1123] = 10'h02B;
    Q_filtered_10b[1122] = 10'h011;
    Q_filtered_10b[1121] = 10'h3F8;
    Q_filtered_10b[1120] = 10'h3DA;
    Q_filtered_10b[1119] = 10'h3B8;
    Q_filtered_10b[1118] = 10'h39D;
    Q_filtered_10b[1117] = 10'h380;
    Q_filtered_10b[1116] = 10'h36B;
    Q_filtered_10b[1115] = 10'h35C;
    Q_filtered_10b[1114] = 10'h356;
    Q_filtered_10b[1113] = 10'h357;
    Q_filtered_10b[1112] = 10'h366;
    Q_filtered_10b[1111] = 10'h381;
    Q_filtered_10b[1110] = 10'h3A2;
    Q_filtered_10b[1109] = 10'h3CE;
    Q_filtered_10b[1108] = 10'h3FB;
    Q_filtered_10b[1107] = 10'h02F;
    Q_filtered_10b[1106] = 10'h062;
    Q_filtered_10b[1105] = 10'h08C;
    Q_filtered_10b[1104] = 10'h0B4;
    Q_filtered_10b[1103] = 10'h0D1;
    Q_filtered_10b[1102] = 10'h0E4;
    Q_filtered_10b[1101] = 10'h0E8;
    Q_filtered_10b[1100] = 10'h0E5;
    Q_filtered_10b[1099] = 10'h0D1;
    Q_filtered_10b[1098] = 10'h0B1;
    Q_filtered_10b[1097] = 10'h086;
    Q_filtered_10b[1096] = 10'h055;
    Q_filtered_10b[1095] = 10'h01F;
    Q_filtered_10b[1094] = 10'h3E4;
    Q_filtered_10b[1093] = 10'h3AB;
    Q_filtered_10b[1092] = 10'h37B;
    Q_filtered_10b[1091] = 10'h34D;
    Q_filtered_10b[1090] = 10'h32C;
    Q_filtered_10b[1089] = 10'h317;
    Q_filtered_10b[1088] = 10'h312;
    Q_filtered_10b[1087] = 10'h315;
    Q_filtered_10b[1086] = 10'h32A;
    Q_filtered_10b[1085] = 10'h34B;
    Q_filtered_10b[1084] = 10'h378;
    Q_filtered_10b[1083] = 10'h3A9;
    Q_filtered_10b[1082] = 10'h3E4;
    Q_filtered_10b[1081] = 10'h023;
    Q_filtered_10b[1080] = 10'h05C;
    Q_filtered_10b[1079] = 10'h090;
    Q_filtered_10b[1078] = 10'h0BA;
    Q_filtered_10b[1077] = 10'h0DB;
    Q_filtered_10b[1076] = 10'h0ED;
    Q_filtered_10b[1075] = 10'h0EE;
    Q_filtered_10b[1074] = 10'h0E4;
    Q_filtered_10b[1073] = 10'h0CC;
    Q_filtered_10b[1072] = 10'h0AB;
    Q_filtered_10b[1071] = 10'h07E;
    Q_filtered_10b[1070] = 10'h050;
    Q_filtered_10b[1069] = 10'h01B;
    Q_filtered_10b[1068] = 10'h3E8;
    Q_filtered_10b[1067] = 10'h3B9;
    Q_filtered_10b[1066] = 10'h38E;
    Q_filtered_10b[1065] = 10'h36A;
    Q_filtered_10b[1064] = 10'h34F;
    Q_filtered_10b[1063] = 10'h33A;
    Q_filtered_10b[1062] = 10'h333;
    Q_filtered_10b[1061] = 10'h32E;
    Q_filtered_10b[1060] = 10'h331;
    Q_filtered_10b[1059] = 10'h33A;
    Q_filtered_10b[1058] = 10'h349;
    Q_filtered_10b[1057] = 10'h353;
    Q_filtered_10b[1056] = 10'h363;
    Q_filtered_10b[1055] = 10'h374;
    Q_filtered_10b[1054] = 10'h37F;
    Q_filtered_10b[1053] = 10'h38B;
    Q_filtered_10b[1052] = 10'h392;
    Q_filtered_10b[1051] = 10'h399;
    Q_filtered_10b[1050] = 10'h39A;
    Q_filtered_10b[1049] = 10'h398;
    Q_filtered_10b[1048] = 10'h394;
    Q_filtered_10b[1047] = 10'h38F;
    Q_filtered_10b[1046] = 10'h388;
    Q_filtered_10b[1045] = 10'h37F;
    Q_filtered_10b[1044] = 10'h377;
    Q_filtered_10b[1043] = 10'h36A;
    Q_filtered_10b[1042] = 10'h35E;
    Q_filtered_10b[1041] = 10'h356;
    Q_filtered_10b[1040] = 10'h34D;
    Q_filtered_10b[1039] = 10'h347;
    Q_filtered_10b[1038] = 10'h342;
    Q_filtered_10b[1037] = 10'h342;
    Q_filtered_10b[1036] = 10'h349;
    Q_filtered_10b[1035] = 10'h351;
    Q_filtered_10b[1034] = 10'h35D;
    Q_filtered_10b[1033] = 10'h368;
    Q_filtered_10b[1032] = 10'h379;
    Q_filtered_10b[1031] = 10'h386;
    Q_filtered_10b[1030] = 10'h398;
    Q_filtered_10b[1029] = 10'h3A5;
    Q_filtered_10b[1028] = 10'h3B1;
    Q_filtered_10b[1027] = 10'h3C1;
    Q_filtered_10b[1026] = 10'h3C9;
    Q_filtered_10b[1025] = 10'h3D2;
    Q_filtered_10b[1024] = 10'h3DB;
    Q_filtered_10b[1023] = 10'h3E4;
    Q_filtered_10b[1022] = 10'h3EB;
    Q_filtered_10b[1021] = 10'h3F7;
    Q_filtered_10b[1020] = 10'h004;
    Q_filtered_10b[1019] = 10'h014;
    Q_filtered_10b[1018] = 10'h02A;
    Q_filtered_10b[1017] = 10'h043;
    Q_filtered_10b[1016] = 10'h05E;
    Q_filtered_10b[1015] = 10'h07B;
    Q_filtered_10b[1014] = 10'h096;
    Q_filtered_10b[1013] = 10'h0AF;
    Q_filtered_10b[1012] = 10'h0C2;
    Q_filtered_10b[1011] = 10'h0CE;
    Q_filtered_10b[1010] = 10'h0D2;
    Q_filtered_10b[1009] = 10'h0CE;
    Q_filtered_10b[1008] = 10'h0BF;
    Q_filtered_10b[1007] = 10'h0A9;
    Q_filtered_10b[1006] = 10'h08E;
    Q_filtered_10b[1005] = 10'h06C;
    Q_filtered_10b[1004] = 10'h049;
    Q_filtered_10b[1003] = 10'h025;
    Q_filtered_10b[1002] = 10'h003;
    Q_filtered_10b[1001] = 10'h3E6;
    Q_filtered_10b[1000] = 10'h3CE;
    Q_filtered_10b[999] = 10'h3BC;
    Q_filtered_10b[998] = 10'h3AD;
    Q_filtered_10b[997] = 10'h3A5;
    Q_filtered_10b[996] = 10'h39F;
    Q_filtered_10b[995] = 10'h39C;
    Q_filtered_10b[994] = 10'h39C;
    Q_filtered_10b[993] = 10'h39E;
    Q_filtered_10b[992] = 10'h39B;
    Q_filtered_10b[991] = 10'h39A;
    Q_filtered_10b[990] = 10'h398;
    Q_filtered_10b[989] = 10'h394;
    Q_filtered_10b[988] = 10'h38F;
    Q_filtered_10b[987] = 10'h38B;
    Q_filtered_10b[986] = 10'h388;
    Q_filtered_10b[985] = 10'h384;
    Q_filtered_10b[984] = 10'h382;
    Q_filtered_10b[983] = 10'h383;
    Q_filtered_10b[982] = 10'h385;
    Q_filtered_10b[981] = 10'h389;
    Q_filtered_10b[980] = 10'h38C;
    Q_filtered_10b[979] = 10'h392;
    Q_filtered_10b[978] = 10'h397;
    Q_filtered_10b[977] = 10'h39B;
    Q_filtered_10b[976] = 10'h39F;
    Q_filtered_10b[975] = 10'h3A3;
    Q_filtered_10b[974] = 10'h3A2;
    Q_filtered_10b[973] = 10'h3A3;
    Q_filtered_10b[972] = 10'h3A6;
    Q_filtered_10b[971] = 10'h3AB;
    Q_filtered_10b[970] = 10'h3B0;
    Q_filtered_10b[969] = 10'h3BC;
    Q_filtered_10b[968] = 10'h3CA;
    Q_filtered_10b[967] = 10'h3DC;
    Q_filtered_10b[966] = 10'h3F4;
    Q_filtered_10b[965] = 10'h00D;
    Q_filtered_10b[964] = 10'h028;
    Q_filtered_10b[963] = 10'h045;
    Q_filtered_10b[962] = 10'h05F;
    Q_filtered_10b[961] = 10'h078;
    Q_filtered_10b[960] = 10'h08B;
    Q_filtered_10b[959] = 10'h099;
    Q_filtered_10b[958] = 10'h09F;
    Q_filtered_10b[957] = 10'h09F;
    Q_filtered_10b[956] = 10'h095;
    Q_filtered_10b[955] = 10'h082;
    Q_filtered_10b[954] = 10'h06B;
    Q_filtered_10b[953] = 10'h04D;
    Q_filtered_10b[952] = 10'h02B;
    Q_filtered_10b[951] = 10'h006;
    Q_filtered_10b[950] = 10'h3E5;
    Q_filtered_10b[949] = 10'h3C7;
    Q_filtered_10b[948] = 10'h3B1;
    Q_filtered_10b[947] = 10'h39F;
    Q_filtered_10b[946] = 10'h395;
    Q_filtered_10b[945] = 10'h395;
    Q_filtered_10b[944] = 10'h39B;
    Q_filtered_10b[943] = 10'h3A6;
    Q_filtered_10b[942] = 10'h3B5;
    Q_filtered_10b[941] = 10'h3CA;
    Q_filtered_10b[940] = 10'h3DE;
    Q_filtered_10b[939] = 10'h3F5;
    Q_filtered_10b[938] = 10'h009;
    Q_filtered_10b[937] = 10'h01A;
    Q_filtered_10b[936] = 10'h02B;
    Q_filtered_10b[935] = 10'h037;
    Q_filtered_10b[934] = 10'h040;
    Q_filtered_10b[933] = 10'h048;
    Q_filtered_10b[932] = 10'h04A;
    Q_filtered_10b[931] = 10'h04F;
    Q_filtered_10b[930] = 10'h054;
    Q_filtered_10b[929] = 10'h05A;
    Q_filtered_10b[928] = 10'h05F;
    Q_filtered_10b[927] = 10'h06B;
    Q_filtered_10b[926] = 10'h077;
    Q_filtered_10b[925] = 10'h085;
    Q_filtered_10b[924] = 10'h094;
    Q_filtered_10b[923] = 10'h0A1;
    Q_filtered_10b[922] = 10'h0AD;
    Q_filtered_10b[921] = 10'h0B6;
    Q_filtered_10b[920] = 10'h0BC;
    Q_filtered_10b[919] = 10'h0BC;
    Q_filtered_10b[918] = 10'h0BA;
    Q_filtered_10b[917] = 10'h0B1;
    Q_filtered_10b[916] = 10'h0A5;
    Q_filtered_10b[915] = 10'h095;
    Q_filtered_10b[914] = 10'h083;
    Q_filtered_10b[913] = 10'h071;
    Q_filtered_10b[912] = 10'h05F;
    Q_filtered_10b[911] = 10'h04D;
    Q_filtered_10b[910] = 10'h03D;
    Q_filtered_10b[909] = 10'h02F;
    Q_filtered_10b[908] = 10'h025;
    Q_filtered_10b[907] = 10'h01A;
    Q_filtered_10b[906] = 10'h011;
    Q_filtered_10b[905] = 10'h00A;
    Q_filtered_10b[904] = 10'h002;
    Q_filtered_10b[903] = 10'h3FD;
    Q_filtered_10b[902] = 10'h3F7;
    Q_filtered_10b[901] = 10'h3F0;
    Q_filtered_10b[900] = 10'h3E6;
    Q_filtered_10b[899] = 10'h3DF;
    Q_filtered_10b[898] = 10'h3D7;
    Q_filtered_10b[897] = 10'h3CC;
    Q_filtered_10b[896] = 10'h3C6;
    Q_filtered_10b[895] = 10'h3C0;
    Q_filtered_10b[894] = 10'h3BA;
    Q_filtered_10b[893] = 10'h3B6;
    Q_filtered_10b[892] = 10'h3B4;
    Q_filtered_10b[891] = 10'h3B1;
    Q_filtered_10b[890] = 10'h3AE;
    Q_filtered_10b[889] = 10'h3AA;
    Q_filtered_10b[888] = 10'h3A4;
    Q_filtered_10b[887] = 10'h39E;
    Q_filtered_10b[886] = 10'h395;
    Q_filtered_10b[885] = 10'h389;
    Q_filtered_10b[884] = 10'h381;
    Q_filtered_10b[883] = 10'h373;
    Q_filtered_10b[882] = 10'h36A;
    Q_filtered_10b[881] = 10'h366;
    Q_filtered_10b[880] = 10'h367;
    Q_filtered_10b[879] = 10'h36B;
    Q_filtered_10b[878] = 10'h37C;
    Q_filtered_10b[877] = 10'h393;
    Q_filtered_10b[876] = 10'h3B1;
    Q_filtered_10b[875] = 10'h3D8;
    Q_filtered_10b[874] = 10'h004;
    Q_filtered_10b[873] = 10'h035;
    Q_filtered_10b[872] = 10'h064;
    Q_filtered_10b[871] = 10'h08E;
    Q_filtered_10b[870] = 10'h0B2;
    Q_filtered_10b[869] = 10'h0CE;
    Q_filtered_10b[868] = 10'h0DF;
    Q_filtered_10b[867] = 10'h0E3;
    Q_filtered_10b[866] = 10'h0DC;
    Q_filtered_10b[865] = 10'h0C9;
    Q_filtered_10b[864] = 10'h0AD;
    Q_filtered_10b[863] = 10'h088;
    Q_filtered_10b[862] = 10'h060;
    Q_filtered_10b[861] = 10'h031;
    Q_filtered_10b[860] = 10'h004;
    Q_filtered_10b[859] = 10'h3DC;
    Q_filtered_10b[858] = 10'h3B7;
    Q_filtered_10b[857] = 10'h39C;
    Q_filtered_10b[856] = 10'h387;
    Q_filtered_10b[855] = 10'h377;
    Q_filtered_10b[854] = 10'h372;
    Q_filtered_10b[853] = 10'h36F;
    Q_filtered_10b[852] = 10'h36E;
    Q_filtered_10b[851] = 10'h36E;
    Q_filtered_10b[850] = 10'h372;
    Q_filtered_10b[849] = 10'h36D;
    Q_filtered_10b[848] = 10'h36A;
    Q_filtered_10b[847] = 10'h363;
    Q_filtered_10b[846] = 10'h358;
    Q_filtered_10b[845] = 10'h350;
    Q_filtered_10b[844] = 10'h347;
    Q_filtered_10b[843] = 10'h340;
    Q_filtered_10b[842] = 10'h33D;
    Q_filtered_10b[841] = 10'h33E;
    Q_filtered_10b[840] = 10'h345;
    Q_filtered_10b[839] = 10'h354;
    Q_filtered_10b[838] = 10'h367;
    Q_filtered_10b[837] = 10'h37E;
    Q_filtered_10b[836] = 10'h39C;
    Q_filtered_10b[835] = 10'h3BA;
    Q_filtered_10b[834] = 10'h3D7;
    Q_filtered_10b[833] = 10'h3F6;
    Q_filtered_10b[832] = 10'h011;
    Q_filtered_10b[831] = 10'h027;
    Q_filtered_10b[830] = 10'h038;
    Q_filtered_10b[829] = 10'h04A;
    Q_filtered_10b[828] = 10'h055;
    Q_filtered_10b[827] = 10'h05F;
    Q_filtered_10b[826] = 10'h068;
    Q_filtered_10b[825] = 10'h06C;
    Q_filtered_10b[824] = 10'h070;
    Q_filtered_10b[823] = 10'h077;
    Q_filtered_10b[822] = 10'h07F;
    Q_filtered_10b[821] = 10'h085;
    Q_filtered_10b[820] = 10'h08E;
    Q_filtered_10b[819] = 10'h098;
    Q_filtered_10b[818] = 10'h0A1;
    Q_filtered_10b[817] = 10'h0A8;
    Q_filtered_10b[816] = 10'h0AE;
    Q_filtered_10b[815] = 10'h0B1;
    Q_filtered_10b[814] = 10'h0B2;
    Q_filtered_10b[813] = 10'h0AF;
    Q_filtered_10b[812] = 10'h0AB;
    Q_filtered_10b[811] = 10'h0A7;
    Q_filtered_10b[810] = 10'h0A1;
    Q_filtered_10b[809] = 10'h09E;
    Q_filtered_10b[808] = 10'h09C;
    Q_filtered_10b[807] = 10'h099;
    Q_filtered_10b[806] = 10'h098;
    Q_filtered_10b[805] = 10'h097;
    Q_filtered_10b[804] = 10'h097;
    Q_filtered_10b[803] = 10'h091;
    Q_filtered_10b[802] = 10'h089;
    Q_filtered_10b[801] = 10'h07E;
    Q_filtered_10b[800] = 10'h06C;
    Q_filtered_10b[799] = 10'h05B;
    Q_filtered_10b[798] = 10'h044;
    Q_filtered_10b[797] = 10'h029;
    Q_filtered_10b[796] = 10'h00D;
    Q_filtered_10b[795] = 10'h3F4;
    Q_filtered_10b[794] = 10'h3D8;
    Q_filtered_10b[793] = 10'h3BE;
    Q_filtered_10b[792] = 10'h3A6;
    Q_filtered_10b[791] = 10'h395;
    Q_filtered_10b[790] = 10'h383;
    Q_filtered_10b[789] = 10'h377;
    Q_filtered_10b[788] = 10'h36E;
    Q_filtered_10b[787] = 10'h368;
    Q_filtered_10b[786] = 10'h367;
    Q_filtered_10b[785] = 10'h367;
    Q_filtered_10b[784] = 10'h366;
    Q_filtered_10b[783] = 10'h366;
    Q_filtered_10b[782] = 10'h369;
    Q_filtered_10b[781] = 10'h367;
    Q_filtered_10b[780] = 10'h366;
    Q_filtered_10b[779] = 10'h360;
    Q_filtered_10b[778] = 10'h35D;
    Q_filtered_10b[777] = 10'h357;
    Q_filtered_10b[776] = 10'h354;
    Q_filtered_10b[775] = 10'h350;
    Q_filtered_10b[774] = 10'h350;
    Q_filtered_10b[773] = 10'h353;
    Q_filtered_10b[772] = 10'h357;
    Q_filtered_10b[771] = 10'h35D;
    Q_filtered_10b[770] = 10'h364;
    Q_filtered_10b[769] = 10'h36D;
    Q_filtered_10b[768] = 10'h376;
    Q_filtered_10b[767] = 10'h37E;
    Q_filtered_10b[766] = 10'h384;
    Q_filtered_10b[765] = 10'h38A;
    Q_filtered_10b[764] = 10'h38E;
    Q_filtered_10b[763] = 10'h393;
    Q_filtered_10b[762] = 10'h393;
    Q_filtered_10b[761] = 10'h394;
    Q_filtered_10b[760] = 10'h391;
    Q_filtered_10b[759] = 10'h390;
    Q_filtered_10b[758] = 10'h38B;
    Q_filtered_10b[757] = 10'h386;
    Q_filtered_10b[756] = 10'h37F;
    Q_filtered_10b[755] = 10'h37C;
    Q_filtered_10b[754] = 10'h379;
    Q_filtered_10b[753] = 10'h379;
    Q_filtered_10b[752] = 10'h378;
    Q_filtered_10b[751] = 10'h37B;
    Q_filtered_10b[750] = 10'h382;
    Q_filtered_10b[749] = 10'h388;
    Q_filtered_10b[748] = 10'h391;
    Q_filtered_10b[747] = 10'h398;
    Q_filtered_10b[746] = 10'h3A2;
    Q_filtered_10b[745] = 10'h3AA;
    Q_filtered_10b[744] = 10'h3B5;
    Q_filtered_10b[743] = 10'h3BB;
    Q_filtered_10b[742] = 10'h3C2;
    Q_filtered_10b[741] = 10'h3CC;
    Q_filtered_10b[740] = 10'h3D1;
    Q_filtered_10b[739] = 10'h3D7;
    Q_filtered_10b[738] = 10'h3DD;
    Q_filtered_10b[737] = 10'h3E4;
    Q_filtered_10b[736] = 10'h3E9;
    Q_filtered_10b[735] = 10'h3F2;
    Q_filtered_10b[734] = 10'h3FC;
    Q_filtered_10b[733] = 10'h009;
    Q_filtered_10b[732] = 10'h019;
    Q_filtered_10b[731] = 10'h02B;
    Q_filtered_10b[730] = 10'h03E;
    Q_filtered_10b[729] = 10'h054;
    Q_filtered_10b[728] = 10'h067;
    Q_filtered_10b[727] = 10'h07B;
    Q_filtered_10b[726] = 10'h08A;
    Q_filtered_10b[725] = 10'h095;
    Q_filtered_10b[724] = 10'h099;
    Q_filtered_10b[723] = 10'h099;
    Q_filtered_10b[722] = 10'h08F;
    Q_filtered_10b[721] = 10'h07D;
    Q_filtered_10b[720] = 10'h067;
    Q_filtered_10b[719] = 10'h04B;
    Q_filtered_10b[718] = 10'h02A;
    Q_filtered_10b[717] = 10'h006;
    Q_filtered_10b[716] = 10'h3E6;
    Q_filtered_10b[715] = 10'h3C8;
    Q_filtered_10b[714] = 10'h3B2;
    Q_filtered_10b[713] = 10'h3A0;
    Q_filtered_10b[712] = 10'h396;
    Q_filtered_10b[711] = 10'h395;
    Q_filtered_10b[710] = 10'h39A;
    Q_filtered_10b[709] = 10'h3A5;
    Q_filtered_10b[708] = 10'h3B4;
    Q_filtered_10b[707] = 10'h3C9;
    Q_filtered_10b[706] = 10'h3DD;
    Q_filtered_10b[705] = 10'h3F5;
    Q_filtered_10b[704] = 10'h00A;
    Q_filtered_10b[703] = 10'h01B;
    Q_filtered_10b[702] = 10'h02D;
    Q_filtered_10b[701] = 10'h038;
    Q_filtered_10b[700] = 10'h041;
    Q_filtered_10b[699] = 10'h048;
    Q_filtered_10b[698] = 10'h04A;
    Q_filtered_10b[697] = 10'h04E;
    Q_filtered_10b[696] = 10'h052;
    Q_filtered_10b[695] = 10'h058;
    Q_filtered_10b[694] = 10'h05D;
    Q_filtered_10b[693] = 10'h06A;
    Q_filtered_10b[692] = 10'h074;
    Q_filtered_10b[691] = 10'h082;
    Q_filtered_10b[690] = 10'h093;
    Q_filtered_10b[689] = 10'h09E;
    Q_filtered_10b[688] = 10'h0AE;
    Q_filtered_10b[687] = 10'h0B8;
    Q_filtered_10b[686] = 10'h0C0;
    Q_filtered_10b[685] = 10'h0C2;
    Q_filtered_10b[684] = 10'h0C2;
    Q_filtered_10b[683] = 10'h0B8;
    Q_filtered_10b[682] = 10'h0A8;
    Q_filtered_10b[681] = 10'h093;
    Q_filtered_10b[680] = 10'h079;
    Q_filtered_10b[679] = 10'h05A;
    Q_filtered_10b[678] = 10'h038;
    Q_filtered_10b[677] = 10'h018;
    Q_filtered_10b[676] = 10'h3FB;
    Q_filtered_10b[675] = 10'h3E4;
    Q_filtered_10b[674] = 10'h3D2;
    Q_filtered_10b[673] = 10'h3C7;
    Q_filtered_10b[672] = 10'h3C3;
    Q_filtered_10b[671] = 10'h3C8;
    Q_filtered_10b[670] = 10'h3D2;
    Q_filtered_10b[669] = 10'h3E1;
    Q_filtered_10b[668] = 10'h3F5;
    Q_filtered_10b[667] = 10'h00B;
    Q_filtered_10b[666] = 10'h023;
    Q_filtered_10b[665] = 10'h03A;
    Q_filtered_10b[664] = 10'h04D;
    Q_filtered_10b[663] = 10'h05E;
    Q_filtered_10b[662] = 10'h06B;
    Q_filtered_10b[661] = 10'h075;
    Q_filtered_10b[660] = 10'h07D;
    Q_filtered_10b[659] = 10'h07E;
    Q_filtered_10b[658] = 10'h082;
    Q_filtered_10b[657] = 10'h084;
    Q_filtered_10b[656] = 10'h086;
    Q_filtered_10b[655] = 10'h086;
    Q_filtered_10b[654] = 10'h08D;
    Q_filtered_10b[653] = 10'h093;
    Q_filtered_10b[652] = 10'h09A;
    Q_filtered_10b[651] = 10'h0A2;
    Q_filtered_10b[650] = 10'h0A8;
    Q_filtered_10b[649] = 10'h0AD;
    Q_filtered_10b[648] = 10'h0B1;
    Q_filtered_10b[647] = 10'h0B3;
    Q_filtered_10b[646] = 10'h0B1;
    Q_filtered_10b[645] = 10'h0AE;
    Q_filtered_10b[644] = 10'h0A7;
    Q_filtered_10b[643] = 10'h0A0;
    Q_filtered_10b[642] = 10'h097;
    Q_filtered_10b[641] = 10'h08D;
    Q_filtered_10b[640] = 10'h084;
    Q_filtered_10b[639] = 10'h07D;
    Q_filtered_10b[638] = 10'h075;
    Q_filtered_10b[637] = 10'h06D;
    Q_filtered_10b[636] = 10'h067;
    Q_filtered_10b[635] = 10'h062;
    Q_filtered_10b[634] = 10'h059;
    Q_filtered_10b[633] = 10'h050;
    Q_filtered_10b[632] = 10'h046;
    Q_filtered_10b[631] = 10'h037;
    Q_filtered_10b[630] = 10'h02A;
    Q_filtered_10b[629] = 10'h019;
    Q_filtered_10b[628] = 10'h005;
    Q_filtered_10b[627] = 10'h3EF;
    Q_filtered_10b[626] = 10'h3DC;
    Q_filtered_10b[625] = 10'h3C6;
    Q_filtered_10b[624] = 10'h3B1;
    Q_filtered_10b[623] = 10'h39D;
    Q_filtered_10b[622] = 10'h38F;
    Q_filtered_10b[621] = 10'h380;
    Q_filtered_10b[620] = 10'h377;
    Q_filtered_10b[619] = 10'h371;
    Q_filtered_10b[618] = 10'h36E;
    Q_filtered_10b[617] = 10'h371;
    Q_filtered_10b[616] = 10'h374;
    Q_filtered_10b[615] = 10'h378;
    Q_filtered_10b[614] = 10'h37C;
    Q_filtered_10b[613] = 10'h382;
    Q_filtered_10b[612] = 10'h385;
    Q_filtered_10b[611] = 10'h387;
    Q_filtered_10b[610] = 10'h387;
    Q_filtered_10b[609] = 10'h388;
    Q_filtered_10b[608] = 10'h387;
    Q_filtered_10b[607] = 10'h388;
    Q_filtered_10b[606] = 10'h388;
    Q_filtered_10b[605] = 10'h38A;
    Q_filtered_10b[604] = 10'h38D;
    Q_filtered_10b[603] = 10'h390;
    Q_filtered_10b[602] = 10'h394;
    Q_filtered_10b[601] = 10'h398;
    Q_filtered_10b[600] = 10'h39B;
    Q_filtered_10b[599] = 10'h3A0;
    Q_filtered_10b[598] = 10'h3A4;
    Q_filtered_10b[597] = 10'h3A7;
    Q_filtered_10b[596] = 10'h3AA;
    Q_filtered_10b[595] = 10'h3AF;
    Q_filtered_10b[594] = 10'h3B6;
    Q_filtered_10b[593] = 10'h3BB;
    Q_filtered_10b[592] = 10'h3C3;
    Q_filtered_10b[591] = 10'h3C9;
    Q_filtered_10b[590] = 10'h3D2;
    Q_filtered_10b[589] = 10'h3DB;
    Q_filtered_10b[588] = 10'h3E7;
    Q_filtered_10b[587] = 10'h3F0;
    Q_filtered_10b[586] = 10'h3FA;
    Q_filtered_10b[585] = 10'h006;
    Q_filtered_10b[584] = 10'h00C;
    Q_filtered_10b[583] = 10'h013;
    Q_filtered_10b[582] = 10'h018;
    Q_filtered_10b[581] = 10'h01C;
    Q_filtered_10b[580] = 10'h01D;
    Q_filtered_10b[579] = 10'h01F;
    Q_filtered_10b[578] = 10'h022;
    Q_filtered_10b[577] = 10'h025;
    Q_filtered_10b[576] = 10'h02B;
    Q_filtered_10b[575] = 10'h032;
    Q_filtered_10b[574] = 10'h03D;
    Q_filtered_10b[573] = 10'h048;
    Q_filtered_10b[572] = 10'h052;
    Q_filtered_10b[571] = 10'h05D;
    Q_filtered_10b[570] = 10'h065;
    Q_filtered_10b[569] = 10'h067;
    Q_filtered_10b[568] = 10'h066;
    Q_filtered_10b[567] = 10'h05E;
    Q_filtered_10b[566] = 10'h04E;
    Q_filtered_10b[565] = 10'h03A;
    Q_filtered_10b[564] = 10'h021;
    Q_filtered_10b[563] = 10'h002;
    Q_filtered_10b[562] = 10'h3E1;
    Q_filtered_10b[561] = 10'h3C0;
    Q_filtered_10b[560] = 10'h39E;
    Q_filtered_10b[559] = 10'h381;
    Q_filtered_10b[558] = 10'h368;
    Q_filtered_10b[557] = 10'h355;
    Q_filtered_10b[556] = 10'h345;
    Q_filtered_10b[555] = 10'h33E;
    Q_filtered_10b[554] = 10'h33A;
    Q_filtered_10b[553] = 10'h33C;
    Q_filtered_10b[552] = 10'h343;
    Q_filtered_10b[551] = 10'h34D;
    Q_filtered_10b[550] = 10'h356;
    Q_filtered_10b[549] = 10'h362;
    Q_filtered_10b[548] = 10'h36F;
    Q_filtered_10b[547] = 10'h378;
    Q_filtered_10b[546] = 10'h381;
    Q_filtered_10b[545] = 10'h385;
    Q_filtered_10b[544] = 10'h38A;
    Q_filtered_10b[543] = 10'h38C;
    Q_filtered_10b[542] = 10'h38D;
    Q_filtered_10b[541] = 10'h38D;
    Q_filtered_10b[540] = 10'h38F;
    Q_filtered_10b[539] = 10'h390;
    Q_filtered_10b[538] = 10'h392;
    Q_filtered_10b[537] = 10'h396;
    Q_filtered_10b[536] = 10'h39A;
    Q_filtered_10b[535] = 10'h39F;
    Q_filtered_10b[534] = 10'h3A5;
    Q_filtered_10b[533] = 10'h3AC;
    Q_filtered_10b[532] = 10'h3AF;
    Q_filtered_10b[531] = 10'h3B3;
    Q_filtered_10b[530] = 10'h3B6;
    Q_filtered_10b[529] = 10'h3BB;
    Q_filtered_10b[528] = 10'h3BC;
    Q_filtered_10b[527] = 10'h3BF;
    Q_filtered_10b[526] = 10'h3C1;
    Q_filtered_10b[525] = 10'h3C6;
    Q_filtered_10b[524] = 10'h3C9;
    Q_filtered_10b[523] = 10'h3D0;
    Q_filtered_10b[522] = 10'h3D8;
    Q_filtered_10b[521] = 10'h3DF;
    Q_filtered_10b[520] = 10'h3E9;
    Q_filtered_10b[519] = 10'h3EF;
    Q_filtered_10b[518] = 10'h3F6;
    Q_filtered_10b[517] = 10'h3F8;
    Q_filtered_10b[516] = 10'h3FA;
    Q_filtered_10b[515] = 10'h3F5;
    Q_filtered_10b[514] = 10'h3EE;
    Q_filtered_10b[513] = 10'h3E5;
    Q_filtered_10b[512] = 10'h3DA;
    Q_filtered_10b[511] = 10'h3CC;
    Q_filtered_10b[510] = 10'h3BC;
    Q_filtered_10b[509] = 10'h3AD;
    Q_filtered_10b[508] = 10'h3A1;
    Q_filtered_10b[507] = 10'h395;
    Q_filtered_10b[506] = 10'h390;
    Q_filtered_10b[505] = 10'h38A;
    Q_filtered_10b[504] = 10'h387;
    Q_filtered_10b[503] = 10'h388;
    Q_filtered_10b[502] = 10'h388;
    Q_filtered_10b[501] = 10'h388;
    Q_filtered_10b[500] = 10'h384;
    Q_filtered_10b[499] = 10'h382;
    Q_filtered_10b[498] = 10'h378;
    Q_filtered_10b[497] = 10'h36F;
    Q_filtered_10b[496] = 10'h360;
    Q_filtered_10b[495] = 10'h351;
    Q_filtered_10b[494] = 10'h346;
    Q_filtered_10b[493] = 10'h339;
    Q_filtered_10b[492] = 10'h330;
    Q_filtered_10b[491] = 10'h32E;
    Q_filtered_10b[490] = 10'h333;
    Q_filtered_10b[489] = 10'h33D;
    Q_filtered_10b[488] = 10'h353;
    Q_filtered_10b[487] = 10'h36E;
    Q_filtered_10b[486] = 10'h391;
    Q_filtered_10b[485] = 10'h3BB;
    Q_filtered_10b[484] = 10'h3EA;
    Q_filtered_10b[483] = 10'h018;
    Q_filtered_10b[482] = 10'h047;
    Q_filtered_10b[481] = 10'h072;
    Q_filtered_10b[480] = 10'h096;
    Q_filtered_10b[479] = 10'h0B2;
    Q_filtered_10b[478] = 10'h0C8;
    Q_filtered_10b[477] = 10'h0D2;
    Q_filtered_10b[476] = 10'h0D5;
    Q_filtered_10b[475] = 10'h0D0;
    Q_filtered_10b[474] = 10'h0C3;
    Q_filtered_10b[473] = 10'h0B2;
    Q_filtered_10b[472] = 10'h0A0;
    Q_filtered_10b[471] = 10'h08C;
    Q_filtered_10b[470] = 10'h077;
    Q_filtered_10b[469] = 10'h068;
    Q_filtered_10b[468] = 10'h05A;
    Q_filtered_10b[467] = 10'h052;
    Q_filtered_10b[466] = 10'h04B;
    Q_filtered_10b[465] = 10'h046;
    Q_filtered_10b[464] = 10'h045;
    Q_filtered_10b[463] = 10'h043;
    Q_filtered_10b[462] = 10'h03E;
    Q_filtered_10b[461] = 10'h039;
    Q_filtered_10b[460] = 10'h035;
    Q_filtered_10b[459] = 10'h02A;
    Q_filtered_10b[458] = 10'h020;
    Q_filtered_10b[457] = 10'h014;
    Q_filtered_10b[456] = 10'h007;
    Q_filtered_10b[455] = 10'h3FB;
    Q_filtered_10b[454] = 10'h3F2;
    Q_filtered_10b[453] = 10'h3EB;
    Q_filtered_10b[452] = 10'h3E4;
    Q_filtered_10b[451] = 10'h3DE;
    Q_filtered_10b[450] = 10'h3DD;
    Q_filtered_10b[449] = 10'h3DC;
    Q_filtered_10b[448] = 10'h3DD;
    Q_filtered_10b[447] = 10'h3DE;
    Q_filtered_10b[446] = 10'h3E1;
    Q_filtered_10b[445] = 10'h3E2;
    Q_filtered_10b[444] = 10'h3E4;
    Q_filtered_10b[443] = 10'h3E4;
    Q_filtered_10b[442] = 10'h3E3;
    Q_filtered_10b[441] = 10'h3E0;
    Q_filtered_10b[440] = 10'h3DF;
    Q_filtered_10b[439] = 10'h3DE;
    Q_filtered_10b[438] = 10'h3DE;
    Q_filtered_10b[437] = 10'h3E1;
    Q_filtered_10b[436] = 10'h3E6;
    Q_filtered_10b[435] = 10'h3EE;
    Q_filtered_10b[434] = 10'h3F7;
    Q_filtered_10b[433] = 10'h004;
    Q_filtered_10b[432] = 10'h010;
    Q_filtered_10b[431] = 10'h01E;
    Q_filtered_10b[430] = 10'h02C;
    Q_filtered_10b[429] = 10'h038;
    Q_filtered_10b[428] = 10'h043;
    Q_filtered_10b[427] = 10'h04B;
    Q_filtered_10b[426] = 10'h052;
    Q_filtered_10b[425] = 10'h055;
    Q_filtered_10b[424] = 10'h057;
    Q_filtered_10b[423] = 10'h055;
    Q_filtered_10b[422] = 10'h050;
    Q_filtered_10b[421] = 10'h049;
    Q_filtered_10b[420] = 10'h041;
    Q_filtered_10b[419] = 10'h039;
    Q_filtered_10b[418] = 10'h02F;
    Q_filtered_10b[417] = 10'h025;
    Q_filtered_10b[416] = 10'h01E;
    Q_filtered_10b[415] = 10'h016;
    Q_filtered_10b[414] = 10'h011;
    Q_filtered_10b[413] = 10'h00D;
    Q_filtered_10b[412] = 10'h00C;
    Q_filtered_10b[411] = 10'h00C;
    Q_filtered_10b[410] = 10'h00E;
    Q_filtered_10b[409] = 10'h014;
    Q_filtered_10b[408] = 10'h01B;
    Q_filtered_10b[407] = 10'h023;
    Q_filtered_10b[406] = 10'h02D;
    Q_filtered_10b[405] = 10'h038;
    Q_filtered_10b[404] = 10'h043;
    Q_filtered_10b[403] = 10'h04B;
    Q_filtered_10b[402] = 10'h054;
    Q_filtered_10b[401] = 10'h05A;
    Q_filtered_10b[400] = 10'h05D;
    Q_filtered_10b[399] = 10'h05B;
    Q_filtered_10b[398] = 10'h057;
    Q_filtered_10b[397] = 10'h04E;
    Q_filtered_10b[396] = 10'h042;
    Q_filtered_10b[395] = 10'h031;
    Q_filtered_10b[394] = 10'h01F;
    Q_filtered_10b[393] = 10'h00A;
    Q_filtered_10b[392] = 10'h3F5;
    Q_filtered_10b[391] = 10'h3E0;
    Q_filtered_10b[390] = 10'h3CD;
    Q_filtered_10b[389] = 10'h3BB;
    Q_filtered_10b[388] = 10'h3AE;
    Q_filtered_10b[387] = 10'h3A4;
    Q_filtered_10b[386] = 10'h3A0;
    Q_filtered_10b[385] = 10'h39F;
    Q_filtered_10b[384] = 10'h3A4;
    Q_filtered_10b[383] = 10'h3AE;
    Q_filtered_10b[382] = 10'h3BB;
    Q_filtered_10b[381] = 10'h3CB;
    Q_filtered_10b[380] = 10'h3DB;
    Q_filtered_10b[379] = 10'h3ED;
    Q_filtered_10b[378] = 10'h3FE;
    Q_filtered_10b[377] = 10'h00C;
    Q_filtered_10b[376] = 10'h01A;
    Q_filtered_10b[375] = 10'h024;
    Q_filtered_10b[374] = 10'h02B;
    Q_filtered_10b[373] = 10'h02D;
    Q_filtered_10b[372] = 10'h02E;
    Q_filtered_10b[371] = 10'h029;
    Q_filtered_10b[370] = 10'h01F;
    Q_filtered_10b[369] = 10'h012;
    Q_filtered_10b[368] = 10'h002;
    Q_filtered_10b[367] = 10'h3EF;
    Q_filtered_10b[366] = 10'h3D8;
    Q_filtered_10b[365] = 10'h3C4;
    Q_filtered_10b[364] = 10'h3B1;
    Q_filtered_10b[363] = 10'h3A2;
    Q_filtered_10b[362] = 10'h396;
    Q_filtered_10b[361] = 10'h392;
    Q_filtered_10b[360] = 10'h395;
    Q_filtered_10b[359] = 10'h39E;
    Q_filtered_10b[358] = 10'h3AF;
    Q_filtered_10b[357] = 10'h3C4;
    Q_filtered_10b[356] = 10'h3E0;
    Q_filtered_10b[355] = 10'h3FF;
    Q_filtered_10b[354] = 10'h023;
    Q_filtered_10b[353] = 10'h045;
    Q_filtered_10b[352] = 10'h066;
    Q_filtered_10b[351] = 10'h085;
    Q_filtered_10b[350] = 10'h09D;
    Q_filtered_10b[349] = 10'h0B0;
    Q_filtered_10b[348] = 10'h0BE;
    Q_filtered_10b[347] = 10'h0C2;
    Q_filtered_10b[346] = 10'h0C3;
    Q_filtered_10b[345] = 10'h0BF;
    Q_filtered_10b[344] = 10'h0B8;
    Q_filtered_10b[343] = 10'h0AD;
    Q_filtered_10b[342] = 10'h0A6;
    Q_filtered_10b[341] = 10'h09D;
    Q_filtered_10b[340] = 10'h098;
    Q_filtered_10b[339] = 10'h094;
    Q_filtered_10b[338] = 10'h090;
    Q_filtered_10b[337] = 10'h08E;
    Q_filtered_10b[336] = 10'h08C;
    Q_filtered_10b[335] = 10'h088;
    Q_filtered_10b[334] = 10'h083;
    Q_filtered_10b[333] = 10'h07B;
    Q_filtered_10b[332] = 10'h06E;
    Q_filtered_10b[331] = 10'h061;
    Q_filtered_10b[330] = 10'h050;
    Q_filtered_10b[329] = 10'h03B;
    Q_filtered_10b[328] = 10'h026;
    Q_filtered_10b[327] = 10'h013;
    Q_filtered_10b[326] = 10'h3FC;
    Q_filtered_10b[325] = 10'h3E9;
    Q_filtered_10b[324] = 10'h3D7;
    Q_filtered_10b[323] = 10'h3CA;
    Q_filtered_10b[322] = 10'h3BB;
    Q_filtered_10b[321] = 10'h3B0;
    Q_filtered_10b[320] = 10'h3A6;
    Q_filtered_10b[319] = 10'h39D;
    Q_filtered_10b[318] = 10'h398;
    Q_filtered_10b[317] = 10'h392;
    Q_filtered_10b[316] = 10'h38A;
    Q_filtered_10b[315] = 10'h383;
    Q_filtered_10b[314] = 10'h37F;
    Q_filtered_10b[313] = 10'h376;
    Q_filtered_10b[312] = 10'h36E;
    Q_filtered_10b[311] = 10'h363;
    Q_filtered_10b[310] = 10'h35C;
    Q_filtered_10b[309] = 10'h353;
    Q_filtered_10b[308] = 10'h34F;
    Q_filtered_10b[307] = 10'h34A;
    Q_filtered_10b[306] = 10'h34A;
    Q_filtered_10b[305] = 10'h34E;
    Q_filtered_10b[304] = 10'h353;
    Q_filtered_10b[303] = 10'h35B;
    Q_filtered_10b[302] = 10'h362;
    Q_filtered_10b[301] = 10'h36C;
    Q_filtered_10b[300] = 10'h376;
    Q_filtered_10b[299] = 10'h37E;
    Q_filtered_10b[298] = 10'h385;
    Q_filtered_10b[297] = 10'h38A;
    Q_filtered_10b[296] = 10'h38E;
    Q_filtered_10b[295] = 10'h393;
    Q_filtered_10b[294] = 10'h393;
    Q_filtered_10b[293] = 10'h394;
    Q_filtered_10b[292] = 10'h392;
    Q_filtered_10b[291] = 10'h390;
    Q_filtered_10b[290] = 10'h38B;
    Q_filtered_10b[289] = 10'h385;
    Q_filtered_10b[288] = 10'h37D;
    Q_filtered_10b[287] = 10'h378;
    Q_filtered_10b[286] = 10'h374;
    Q_filtered_10b[285] = 10'h373;
    Q_filtered_10b[284] = 10'h371;
    Q_filtered_10b[283] = 10'h375;
    Q_filtered_10b[282] = 10'h37D;
    Q_filtered_10b[281] = 10'h385;
    Q_filtered_10b[280] = 10'h392;
    Q_filtered_10b[279] = 10'h39C;
    Q_filtered_10b[278] = 10'h3AC;
    Q_filtered_10b[277] = 10'h3B9;
    Q_filtered_10b[276] = 10'h3CB;
    Q_filtered_10b[275] = 10'h3D8;
    Q_filtered_10b[274] = 10'h3E5;
    Q_filtered_10b[273] = 10'h3F5;
    Q_filtered_10b[272] = 10'h3FE;
    Q_filtered_10b[271] = 10'h007;
    Q_filtered_10b[270] = 10'h010;
    Q_filtered_10b[269] = 10'h017;
    Q_filtered_10b[268] = 10'h01C;
    Q_filtered_10b[267] = 10'h025;
    Q_filtered_10b[266] = 10'h02E;
    Q_filtered_10b[265] = 10'h03A;
    Q_filtered_10b[264] = 10'h04B;
    Q_filtered_10b[263] = 10'h05E;
    Q_filtered_10b[262] = 10'h074;
    Q_filtered_10b[261] = 10'h08C;
    Q_filtered_10b[260] = 10'h0A2;
    Q_filtered_10b[259] = 10'h0B7;
    Q_filtered_10b[258] = 10'h0C7;
    Q_filtered_10b[257] = 10'h0D1;
    Q_filtered_10b[256] = 10'h0D2;
    Q_filtered_10b[255] = 10'h0CC;
    Q_filtered_10b[254] = 10'h0BB;
    Q_filtered_10b[253] = 10'h0A2;
    Q_filtered_10b[252] = 10'h082;
    Q_filtered_10b[251] = 10'h05B;
    Q_filtered_10b[250] = 10'h032;
    Q_filtered_10b[249] = 10'h008;
    Q_filtered_10b[248] = 10'h3DE;
    Q_filtered_10b[247] = 10'h3BA;
    Q_filtered_10b[246] = 10'h39B;
    Q_filtered_10b[245] = 10'h383;
    Q_filtered_10b[244] = 10'h370;
    Q_filtered_10b[243] = 10'h367;
    Q_filtered_10b[242] = 10'h361;
    Q_filtered_10b[241] = 10'h363;
    Q_filtered_10b[240] = 10'h36B;
    Q_filtered_10b[239] = 10'h378;
    Q_filtered_10b[238] = 10'h383;
    Q_filtered_10b[237] = 10'h392;
    Q_filtered_10b[236] = 10'h3A3;
    Q_filtered_10b[235] = 10'h3AF;
    Q_filtered_10b[234] = 10'h3BA;
    Q_filtered_10b[233] = 10'h3C1;
    Q_filtered_10b[232] = 10'h3C7;
    Q_filtered_10b[231] = 10'h3C8;
    Q_filtered_10b[230] = 10'h3C6;
    Q_filtered_10b[229] = 10'h3C2;
    Q_filtered_10b[228] = 10'h3BD;
    Q_filtered_10b[227] = 10'h3B7;
    Q_filtered_10b[226] = 10'h3AE;
    Q_filtered_10b[225] = 10'h3A7;
    Q_filtered_10b[224] = 10'h39E;
    Q_filtered_10b[223] = 10'h395;
    Q_filtered_10b[222] = 10'h38E;
    Q_filtered_10b[221] = 10'h387;
    Q_filtered_10b[220] = 10'h380;
    Q_filtered_10b[219] = 10'h37C;
    Q_filtered_10b[218] = 10'h37A;
    Q_filtered_10b[217] = 10'h37D;
    Q_filtered_10b[216] = 10'h37F;
    Q_filtered_10b[215] = 10'h386;
    Q_filtered_10b[214] = 10'h38D;
    Q_filtered_10b[213] = 10'h399;
    Q_filtered_10b[212] = 10'h3A3;
    Q_filtered_10b[211] = 10'h3B1;
    Q_filtered_10b[210] = 10'h3BD;
    Q_filtered_10b[209] = 10'h3CA;
    Q_filtered_10b[208] = 10'h3D7;
    Q_filtered_10b[207] = 10'h3E1;
    Q_filtered_10b[206] = 10'h3E9;
    Q_filtered_10b[205] = 10'h3F0;
    Q_filtered_10b[204] = 10'h3F4;
    Q_filtered_10b[203] = 10'h3F5;
    Q_filtered_10b[202] = 10'h3F6;
    Q_filtered_10b[201] = 10'h3F3;
    Q_filtered_10b[200] = 10'h3F1;
    Q_filtered_10b[199] = 10'h3EE;
    Q_filtered_10b[198] = 10'h3EB;
    Q_filtered_10b[197] = 10'h3E8;
    Q_filtered_10b[196] = 10'h3E7;
    Q_filtered_10b[195] = 10'h3E7;
    Q_filtered_10b[194] = 10'h3E6;
    Q_filtered_10b[193] = 10'h3E7;
    Q_filtered_10b[192] = 10'h3E7;
    Q_filtered_10b[191] = 10'h3E9;
    Q_filtered_10b[190] = 10'h3E9;
    Q_filtered_10b[189] = 10'h3E9;
    Q_filtered_10b[188] = 10'h3E9;
    Q_filtered_10b[187] = 10'h3EA;
    Q_filtered_10b[186] = 10'h3E9;
    Q_filtered_10b[185] = 10'h3EA;
    Q_filtered_10b[184] = 10'h3EB;
    Q_filtered_10b[183] = 10'h3EB;
    Q_filtered_10b[182] = 10'h3ED;
    Q_filtered_10b[181] = 10'h3EE;
    Q_filtered_10b[180] = 10'h3F0;
    Q_filtered_10b[179] = 10'h3EF;
    Q_filtered_10b[178] = 10'h3EF;
    Q_filtered_10b[177] = 10'h3EC;
    Q_filtered_10b[176] = 10'h3E8;
    Q_filtered_10b[175] = 10'h3E4;
    Q_filtered_10b[174] = 10'h3DF;
    Q_filtered_10b[173] = 10'h3D8;
    Q_filtered_10b[172] = 10'h3D3;
    Q_filtered_10b[171] = 10'h3CE;
    Q_filtered_10b[170] = 10'h3C8;
    Q_filtered_10b[169] = 10'h3C4;
    Q_filtered_10b[168] = 10'h3BE;
    Q_filtered_10b[167] = 10'h3BB;
    Q_filtered_10b[166] = 10'h3B7;
    Q_filtered_10b[165] = 10'h3B6;
    Q_filtered_10b[164] = 10'h3B2;
    Q_filtered_10b[163] = 10'h3B1;
    Q_filtered_10b[162] = 10'h3B1;
    Q_filtered_10b[161] = 10'h3B2;
    Q_filtered_10b[160] = 10'h3B3;
    Q_filtered_10b[159] = 10'h3B5;
    Q_filtered_10b[158] = 10'h3B9;
    Q_filtered_10b[157] = 10'h3BC;
    Q_filtered_10b[156] = 10'h3BF;
    Q_filtered_10b[155] = 10'h3C0;
    Q_filtered_10b[154] = 10'h3C2;
    Q_filtered_10b[153] = 10'h3C1;
    Q_filtered_10b[152] = 10'h3C1;
    Q_filtered_10b[151] = 10'h3BC;
    Q_filtered_10b[150] = 10'h3B8;
    Q_filtered_10b[149] = 10'h3B3;
    Q_filtered_10b[148] = 10'h3AE;
    Q_filtered_10b[147] = 10'h3A7;
    Q_filtered_10b[146] = 10'h39F;
    Q_filtered_10b[145] = 10'h398;
    Q_filtered_10b[144] = 10'h392;
    Q_filtered_10b[143] = 10'h38D;
    Q_filtered_10b[142] = 10'h38A;
    Q_filtered_10b[141] = 10'h387;
    Q_filtered_10b[140] = 10'h386;
    Q_filtered_10b[139] = 10'h388;
    Q_filtered_10b[138] = 10'h388;
    Q_filtered_10b[137] = 10'h38A;
    Q_filtered_10b[136] = 10'h389;
    Q_filtered_10b[135] = 10'h38A;
    Q_filtered_10b[134] = 10'h387;
    Q_filtered_10b[133] = 10'h385;
    Q_filtered_10b[132] = 10'h37F;
    Q_filtered_10b[131] = 10'h37A;
    Q_filtered_10b[130] = 10'h377;
    Q_filtered_10b[129] = 10'h373;
    Q_filtered_10b[128] = 10'h370;
    Q_filtered_10b[127] = 10'h372;
    Q_filtered_10b[126] = 10'h377;
    Q_filtered_10b[125] = 10'h37E;
    Q_filtered_10b[124] = 10'h38C;
    Q_filtered_10b[123] = 10'h39A;
    Q_filtered_10b[122] = 10'h3AE;
    Q_filtered_10b[121] = 10'h3C4;
    Q_filtered_10b[120] = 10'h3DE;
    Q_filtered_10b[119] = 10'h3F6;
    Q_filtered_10b[118] = 10'h00F;
    Q_filtered_10b[117] = 10'h027;
    Q_filtered_10b[116] = 10'h039;
    Q_filtered_10b[115] = 10'h048;
    Q_filtered_10b[114] = 10'h054;
    Q_filtered_10b[113] = 10'h05B;
    Q_filtered_10b[112] = 10'h05C;
    Q_filtered_10b[111] = 10'h05C;
    Q_filtered_10b[110] = 10'h059;
    Q_filtered_10b[109] = 10'h055;
    Q_filtered_10b[108] = 10'h053;
    Q_filtered_10b[107] = 10'h050;
    Q_filtered_10b[106] = 10'h04F;
    Q_filtered_10b[105] = 10'h051;
    Q_filtered_10b[104] = 10'h052;
    Q_filtered_10b[103] = 10'h057;
    Q_filtered_10b[102] = 10'h05A;
    Q_filtered_10b[101] = 10'h05B;
    Q_filtered_10b[100] = 10'h05B;
    Q_filtered_10b[99] = 10'h056;
    Q_filtered_10b[98] = 10'h04B;
    Q_filtered_10b[97] = 10'h03C;
    Q_filtered_10b[96] = 10'h02A;
    Q_filtered_10b[95] = 10'h011;
    Q_filtered_10b[94] = 10'h3F5;
    Q_filtered_10b[93] = 10'h3D8;
    Q_filtered_10b[92] = 10'h3BB;
    Q_filtered_10b[91] = 10'h3A1;
    Q_filtered_10b[90] = 10'h38C;
    Q_filtered_10b[89] = 10'h37C;
    Q_filtered_10b[88] = 10'h370;
    Q_filtered_10b[87] = 10'h36C;
    Q_filtered_10b[86] = 10'h36E;
    Q_filtered_10b[85] = 10'h374;
    Q_filtered_10b[84] = 10'h37F;
    Q_filtered_10b[83] = 10'h38D;
    Q_filtered_10b[82] = 10'h39B;
    Q_filtered_10b[81] = 10'h3AA;
    Q_filtered_10b[80] = 10'h3B7;
    Q_filtered_10b[79] = 10'h3C2;
    Q_filtered_10b[78] = 10'h3CC;
    Q_filtered_10b[77] = 10'h3D3;
    Q_filtered_10b[76] = 10'h3D9;
    Q_filtered_10b[75] = 10'h3DF;
    Q_filtered_10b[74] = 10'h3E4;
    Q_filtered_10b[73] = 10'h3EB;
    Q_filtered_10b[72] = 10'h3F4;
    Q_filtered_10b[71] = 10'h3FE;
    Q_filtered_10b[70] = 10'h009;
    Q_filtered_10b[69] = 10'h019;
    Q_filtered_10b[68] = 10'h02A;
    Q_filtered_10b[67] = 10'h03A;
    Q_filtered_10b[66] = 10'h04C;
    Q_filtered_10b[65] = 10'h05C;
    Q_filtered_10b[64] = 10'h069;
    Q_filtered_10b[63] = 10'h074;
    Q_filtered_10b[62] = 10'h07E;
    Q_filtered_10b[61] = 10'h083;
    Q_filtered_10b[60] = 10'h087;
    Q_filtered_10b[59] = 10'h088;
    Q_filtered_10b[58] = 10'h086;
    Q_filtered_10b[57] = 10'h084;
    Q_filtered_10b[56] = 10'h083;
    Q_filtered_10b[55] = 10'h081;
    Q_filtered_10b[54] = 10'h080;
    Q_filtered_10b[53] = 10'h080;
    Q_filtered_10b[52] = 10'h080;
    Q_filtered_10b[51] = 10'h084;
    Q_filtered_10b[50] = 10'h085;
    Q_filtered_10b[49] = 10'h086;
    Q_filtered_10b[48] = 10'h083;
    Q_filtered_10b[47] = 10'h080;
    Q_filtered_10b[46] = 10'h078;
    Q_filtered_10b[45] = 10'h06D;
    Q_filtered_10b[44] = 10'h05F;
    Q_filtered_10b[43] = 10'h04E;
    Q_filtered_10b[42] = 10'h03C;
    Q_filtered_10b[41] = 10'h029;
    Q_filtered_10b[40] = 10'h014;
    Q_filtered_10b[39] = 10'h002;
    Q_filtered_10b[38] = 10'h3F3;
    Q_filtered_10b[37] = 10'h3E7;
    Q_filtered_10b[36] = 10'h3DC;
    Q_filtered_10b[35] = 10'h3D6;
    Q_filtered_10b[34] = 10'h3D4;
    Q_filtered_10b[33] = 10'h3D4;
    Q_filtered_10b[32] = 10'h3D9;
    Q_filtered_10b[31] = 10'h3DE;
    Q_filtered_10b[30] = 10'h3E5;
    Q_filtered_10b[29] = 10'h3ED;
    Q_filtered_10b[28] = 10'h3F5;
    Q_filtered_10b[27] = 10'h3FB;
    Q_filtered_10b[26] = 10'h000;
    Q_filtered_10b[25] = 10'h002;
    Q_filtered_10b[24] = 10'h004;
    Q_filtered_10b[23] = 10'h004;
    Q_filtered_10b[22] = 10'h003;
    Q_filtered_10b[21] = 10'h002;
    Q_filtered_10b[20] = 10'h000;
    Q_filtered_10b[19] = 10'h000;
    Q_filtered_10b[18] = 10'h3FE;
    Q_filtered_10b[17] = 10'h3FF;
    Q_filtered_10b[16] = 10'h3FE;
    Q_filtered_10b[15] = 10'h3FF;
    Q_filtered_10b[14] = 10'h000;
    Q_filtered_10b[13] = 10'h3FF;
    Q_filtered_10b[12] = 10'h3FF;
    Q_filtered_10b[11] = 10'h3FF;
    Q_filtered_10b[10] = 10'h000;
    Q_filtered_10b[9] = 10'h000;
    Q_filtered_10b[8] = 10'h000;
    Q_filtered_10b[7] = 10'h000;
    Q_filtered_10b[6] = 10'h000;
    Q_filtered_10b[5] = 10'h001;
    Q_filtered_10b[4] = 10'h000;
    Q_filtered_10b[3] = 10'h000;
    Q_filtered_10b[2] = 10'h000;
    Q_filtered_10b[1] = 10'h000;
    Q_filtered_10b[0] = 10'h000;


// I Channel 12b Expected output
//     first 64 samples only
    I_filtered_12b[63] = 12'h000;
    I_filtered_12b[62] = 12'h000;
    I_filtered_12b[61] = 12'h005;
    I_filtered_12b[60] = 12'h00A;
    I_filtered_12b[59] = 12'h00A;
    I_filtered_12b[58] = 12'h00F;
    I_filtered_12b[57] = 12'h00A;
    I_filtered_12b[56] = 12'h00A;
    I_filtered_12b[55] = 12'h005;
    I_filtered_12b[54] = 12'h000;
    I_filtered_12b[53] = 12'hFF6;
    I_filtered_12b[52] = 12'hFF1;
    I_filtered_12b[51] = 12'hFF1;
    I_filtered_12b[50] = 12'hFF1;
    I_filtered_12b[49] = 12'hFF6;
    I_filtered_12b[48] = 12'hFFA;
    I_filtered_12b[47] = 12'h008;
    I_filtered_12b[46] = 12'h017;
    I_filtered_12b[45] = 12'h025;
    I_filtered_12b[44] = 12'h035;
    I_filtered_12b[43] = 12'h03F;
    I_filtered_12b[42] = 12'h040;
    I_filtered_12b[41] = 12'h03C;
    I_filtered_12b[40] = 12'h02F;
    I_filtered_12b[39] = 12'h00D;
    I_filtered_12b[38] = 12'hFE0;
    I_filtered_12b[37] = 12'hFA9;
    I_filtered_12b[36] = 12'hF62;
    I_filtered_12b[35] = 12'hF10;
    I_filtered_12b[34] = 12'hEBC;
    I_filtered_12b[33] = 12'hE64;
    I_filtered_12b[32] = 12'hE15;
    I_filtered_12b[31] = 12'hDD2;
    I_filtered_12b[30] = 12'hD9E;
    I_filtered_12b[29] = 12'hD81;
    I_filtered_12b[28] = 12'hD79;
    I_filtered_12b[27] = 12'hD88;
    I_filtered_12b[26] = 12'hDAE;
    I_filtered_12b[25] = 12'hDE9;
    I_filtered_12b[24] = 12'hE35;
    I_filtered_12b[23] = 12'hE8D;
    I_filtered_12b[22] = 12'hEEE;
    I_filtered_12b[21] = 12'hF48;
    I_filtered_12b[20] = 12'hFA6;
    I_filtered_12b[19] = 12'hFF5;
    I_filtered_12b[18] = 12'h039;
    I_filtered_12b[17] = 12'h06E;
    I_filtered_12b[16] = 12'h09A;
    I_filtered_12b[15] = 12'h0AF;
    I_filtered_12b[14] = 12'h0BB;
    I_filtered_12b[13] = 12'h0BF;
    I_filtered_12b[12] = 12'h0B4;
    I_filtered_12b[11] = 12'h0A3;
    I_filtered_12b[10] = 12'h090;
    I_filtered_12b[9] = 12'h082;
    I_filtered_12b[8] = 12'h06F;
    I_filtered_12b[7] = 12'h062;
    I_filtered_12b[6] = 12'h05A;
    I_filtered_12b[5] = 12'h04E;
    I_filtered_12b[4] = 12'h049;
    I_filtered_12b[3] = 12'h048;
    I_filtered_12b[2] = 12'h04F;
    I_filtered_12b[1] = 12'h050;
    I_filtered_12b[0] = 12'h05F;


// Q Channel 12b Expected output
//     first 64 samples only
    Q_filtered_12b[63] = 12'h000;
    Q_filtered_12b[62] = 12'h000;
    Q_filtered_12b[61] = 12'h001;
    Q_filtered_12b[60] = 12'h002;
    Q_filtered_12b[59] = 12'h002;
    Q_filtered_12b[58] = 12'h003;
    Q_filtered_12b[57] = 12'h002;
    Q_filtered_12b[56] = 12'h002;
    Q_filtered_12b[55] = 12'h001;
    Q_filtered_12b[54] = 12'h000;
    Q_filtered_12b[53] = 12'hFFE;
    Q_filtered_12b[52] = 12'hFFD;
    Q_filtered_12b[51] = 12'hFFD;
    Q_filtered_12b[50] = 12'hFFD;
    Q_filtered_12b[49] = 12'hFFE;
    Q_filtered_12b[48] = 12'hFFA;
    Q_filtered_12b[47] = 12'hFF8;
    Q_filtered_12b[46] = 12'hFFB;
    Q_filtered_12b[45] = 12'hFF8;
    Q_filtered_12b[44] = 12'h000;
    Q_filtered_12b[43] = 12'h002;
    Q_filtered_12b[42] = 12'h007;
    Q_filtered_12b[41] = 12'h00B;
    Q_filtered_12b[40] = 12'h012;
    Q_filtered_12b[39] = 12'h011;
    Q_filtered_12b[38] = 12'h009;
    Q_filtered_12b[37] = 12'hFFF;
    Q_filtered_12b[36] = 12'hFED;
    Q_filtered_12b[35] = 12'hFD5;
    Q_filtered_12b[34] = 12'hFB2;
    Q_filtered_12b[33] = 12'hF94;
    Q_filtered_12b[32] = 12'hF78;
    Q_filtered_12b[31] = 12'hF62;
    Q_filtered_12b[30] = 12'hF4F;
    Q_filtered_12b[29] = 12'hF4E;
    Q_filtered_12b[28] = 12'hF57;
    Q_filtered_12b[27] = 12'hF71;
    Q_filtered_12b[26] = 12'hF9A;
    Q_filtered_12b[25] = 12'hFCB;
    Q_filtered_12b[24] = 12'h009;
    Q_filtered_12b[23] = 12'h052;
    Q_filtered_12b[22] = 12'h0A3;
    Q_filtered_12b[21] = 12'h0EF;
    Q_filtered_12b[20] = 12'h139;
    Q_filtered_12b[19] = 12'h17E;
    Q_filtered_12b[18] = 12'h1B4;
    Q_filtered_12b[17] = 12'h1DF;
    Q_filtered_12b[16] = 12'h202;
    Q_filtered_12b[15] = 12'h20E;
    Q_filtered_12b[14] = 12'h217;
    Q_filtered_12b[13] = 12'h216;
    Q_filtered_12b[12] = 12'h20F;
    Q_filtered_12b[11] = 12'h202;
    Q_filtered_12b[10] = 12'h201;
    Q_filtered_12b[9] = 12'h1FF;
    Q_filtered_12b[8] = 12'h204;
    Q_filtered_12b[7] = 12'h20B;
    Q_filtered_12b[6] = 12'h211;
    Q_filtered_12b[5] = 12'h219;
    Q_filtered_12b[4] = 12'h220;
    Q_filtered_12b[3] = 12'h21C;
    Q_filtered_12b[2] = 12'h20E;
    Q_filtered_12b[1] = 12'h1F8;
    Q_filtered_12b[0] = 12'h1D0;
end

endmodule

