`timescale 1ns / 1ps
`include "modulator_signals.vh"

module baseband_dsp_tb;

    reg data_in;
    reg data_clk;
    reg dsp_clk;
    reg rst_n_data;
    reg rst_n_dsp;
    reg msg_in;
    reg rw;
    reg [9:0] mem_addr;
    reg [7:0] coeff_in;
    reg enable;
    reg [3:0] sample_rate;
    reg mapping;
    wire mem_read_out;
    wire [9:0] I_out;
    wire [9:0] Q_out; 

    baseband_dsp DUT(
        .data_in(data_in),
        .data_clk(data_clk),
        .dsp_clk(dsp_clk),
        .rst_n_data(rst_n_data),
        .rst_n_dsp(rst_n_dsp),
        .msg_in(msg_in),
        .rw(rw),
        .mem_addr(mem_addr),
        .coeff_in(coeff_in),
        .mem_read_out(mem_read_out),
        .I_out(I_out),
	    .Q_out(Q_out)
    );
	
	// Datastream variables
	reg [7:0] Icoeff [0:70];
	reg [7:0] Qcoeff [0:70];	
	reg [779:0] datastream;
	reg [9:0] I_filtered_10b[0:1733];
	reg [9:0] Q_filtered_10b[0:1733];
	reg [11:0] I_filtered_12b[0:63];
	reg [11:0] Q_filtered_12b[0:63];
	
    always #8.333 data_clk = ~data_clk;
    always #3.846 dsp_clk = ~dsp_clk;
    
    reg [8*39:0] testcase;
    integer i;
	
    initial begin
        testcase = "Initializing";
        data_clk <= 1'b0;
        dsp_clk <= 1'b0;
        rst_n_data <= 1'b0;
        rst_n_dsp <= 1'b0;
		sample_rate <= 4'd13;
        data_in <= 1'b0; 
        enable <= 1'b0;

		repeat(2) @(posedge data_clk);
		rst_n_data <= 1'b1;
        enable <= 1'b1;
		@(posedge data_clk);

        @(posedge dsp_clk)
        rst_n_dsp <= 1'b1;
        @(posedge dsp_clk)

        // Write I coefficients to memory
        @(negedge dsp_clk);
		for (i=0; i<=70; i=i+1) begin
			msg_in <= 1'b1;
			rw <= 1'b1;
			mem_addr  <= i + 128;
			coeff_in  <= Icoeff[i];
			@(negedge dsp_clk);	 
		end

		// Write Q coefficients to memory
		for (i=0; i<=70; i = i+1) begin
			msg_in <= 1'b1;
			rw <= 1'b1;
			mem_addr  <= i + 256;
			coeff_in  <= Qcoeff[i];
			@(negedge dsp_clk);	 
		end
		msg_in <= 1'b0;

        testcase = "Coeff_Read";
        repeat(3) @(posedge dsp_clk);
        // Test reading coeff I memory
		// coeff_read_out should set to 0xFD
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr  <= 133; // This is addr of 5th I coeff: oxFD
		repeat(2) @(posedge dsp_clk);
		msg_in <= 1'b0;

		repeat(3) @(posedge dsp_clk);
		// Test reading coeff Q memory
		// coeff_read_out should set to 0x02
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr  <= 266; 
		repeat(3) @(posedge dsp_clk);
		msg_in <= 1'b0;

		// flush the pipeline
		repeat(5) @(posedge dsp_clk);

        // Send in datastream with 12 bit header
        testcase <= "Datastream";    
        @(negedge data_clk);
        for (i=779; i>=0; i=i-1) begin
            data_in <= datastream[i]; 
            @(negedge data_clk);
        end

        repeat(3) @(posedge dsp_clk);
        // Test reading I output memory
		// Should read 10th output: 0x00 or 0x05F idk
        testcase <= "Output_read"; 
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr <= 512;
		// Read last 4 LSBs
		repeat(1) @(posedge dsp_clk);
		mem_addr  <= 513;
		repeat(3) @(posedge dsp_clk);

		// Test reading I output memory
		// Should read 10th output: 0x090 or 0x082 or 0xFF6 idk
        testcase <= "Output_read"; 
		msg_in <= 1'b1;
		rw <= 1'b0;
		mem_addr <= 532;
		// Read last 4 LSBs
		repeat(1) @(posedge dsp_clk);
		mem_addr  <= 533;
		repeat(3) @(posedge dsp_clk);

        // Write compare outputs function and log file
        $finish;
    end

initial begin
    // I filter coefficients
    reg [7:0] Icoeff[0] = 00;
    reg [7:0] Icoeff[1] = 00;
    reg [7:0] Icoeff[2] = FF;
    reg [7:0] Icoeff[3] = FE;
    reg [7:0] Icoeff[4] = FE;
    reg [7:0] Icoeff[5] = FD;
    reg [7:0] Icoeff[6] = FE;
    reg [7:0] Icoeff[7] = FE;
    reg [7:0] Icoeff[8] = FF;
    reg [7:0] Icoeff[9] = 00;
    reg [7:0] Icoeff[10] = 02;
    reg [7:0] Icoeff[11] = 03;
    reg [7:0] Icoeff[12] = 03;
    reg [7:0] Icoeff[13] = 03;
    reg [7:0] Icoeff[14] = 02;
    reg [7:0] Icoeff[15] = 01;
    reg [7:0] Icoeff[16] = FE;
    reg [7:0] Icoeff[17] = FB;
    reg [7:0] Icoeff[18] = F8;
    reg [7:0] Icoeff[19] = F5;
    reg [7:0] Icoeff[20] = F3;
    reg [7:0] Icoeff[21] = F3;
    reg [7:0] Icoeff[22] = F4;
    reg [7:0] Icoeff[23] = F7;
    reg [7:0] Icoeff[24] = FE;
    reg [7:0] Icoeff[25] = 07;
    reg [7:0] Icoeff[26] = 12;
    reg [7:0] Icoeff[27] = 20;
    reg [7:0] Icoeff[28] = 30;
    reg [7:0] Icoeff[29] = 40;
    reg [7:0] Icoeff[30] = 51;
    reg [7:0] Icoeff[31] = 60;
    reg [7:0] Icoeff[32] = 6D;
    reg [7:0] Icoeff[33] = 77;
    reg [7:0] Icoeff[34] = 7D;
    reg [7:0] Icoeff[35] = 7F;
    reg [7:0] Icoeff[36] = 7D;
    reg [7:0] Icoeff[37] = 77;
    reg [7:0] Icoeff[38] = 6D;
    reg [7:0] Icoeff[39] = 60;
    reg [7:0] Icoeff[40] = 51;
    reg [7:0] Icoeff[41] = 40;
    reg [7:0] Icoeff[42] = 30;
    reg [7:0] Icoeff[43] = 20;
    reg [7:0] Icoeff[44] = 12;
    reg [7:0] Icoeff[45] = 07;
    reg [7:0] Icoeff[46] = FE;
    reg [7:0] Icoeff[47] = F7;
    reg [7:0] Icoeff[48] = F4;
    reg [7:0] Icoeff[49] = F3;
    reg [7:0] Icoeff[50] = F3;
    reg [7:0] Icoeff[51] = F5;
    reg [7:0] Icoeff[52] = F8;
    reg [7:0] Icoeff[53] = FB;
    reg [7:0] Icoeff[54] = FE;
    reg [7:0] Icoeff[55] = 01;
    reg [7:0] Icoeff[56] = 02;
    reg [7:0] Icoeff[57] = 03;
    reg [7:0] Icoeff[58] = 03;
    reg [7:0] Icoeff[59] = 03;
    reg [7:0] Icoeff[60] = 02;
    reg [7:0] Icoeff[61] = 00;
    reg [7:0] Icoeff[62] = FF;
    reg [7:0] Icoeff[63] = FE;
    reg [7:0] Icoeff[64] = FE;
    reg [7:0] Icoeff[65] = FD;
    reg [7:0] Icoeff[66] = FE;
    reg [7:0] Icoeff[67] = FE;
    reg [7:0] Icoeff[68] = FF;
    reg [7:0] Icoeff[69] = 00;
    reg [7:0] Icoeff[70] = 00;


    // Q filter coefficients
    reg [7:0] Qcoeff[0] = 00;
    reg [7:0] Qcoeff[1] = 00;
    reg [7:0] Qcoeff[2] = FF;
    reg [7:0] Qcoeff[3] = FE;
    reg [7:0] Qcoeff[4] = FE;
    reg [7:0] Qcoeff[5] = FD;
    reg [7:0] Qcoeff[6] = FE;
    reg [7:0] Qcoeff[7] = FE;
    reg [7:0] Qcoeff[8] = FF;
    reg [7:0] Qcoeff[9] = 00;
    reg [7:0] Qcoeff[10] = 02;
    reg [7:0] Qcoeff[11] = 03;
    reg [7:0] Qcoeff[12] = 03;
    reg [7:0] Qcoeff[13] = 03;
    reg [7:0] Qcoeff[14] = 02;
    reg [7:0] Qcoeff[15] = 01;
    reg [7:0] Qcoeff[16] = FE;
    reg [7:0] Qcoeff[17] = FB;
    reg [7:0] Qcoeff[18] = F9;
    reg [7:0] Qcoeff[19] = F6;
    reg [7:0] Qcoeff[20] = F4;
    reg [7:0] Qcoeff[21] = F4;
    reg [7:0] Qcoeff[22] = F5;
    reg [7:0] Qcoeff[23] = F8;
    reg [7:0] Qcoeff[24] = FE;
    reg [7:0] Qcoeff[25] = 06;
    reg [7:0] Qcoeff[26] = 10;
    reg [7:0] Qcoeff[27] = 1D;
    reg [7:0] Qcoeff[28] = 2B;
    reg [7:0] Qcoeff[29] = 3A;
    reg [7:0] Qcoeff[30] = 49;
    reg [7:0] Qcoeff[31] = 56;
    reg [7:0] Qcoeff[32] = 62;
    reg [7:0] Qcoeff[33] = 6B;
    reg [7:0] Qcoeff[34] = 71;
    reg [7:0] Qcoeff[35] = 72;
    reg [7:0] Qcoeff[36] = 71;
    reg [7:0] Qcoeff[37] = 6B;
    reg [7:0] Qcoeff[38] = 62;
    reg [7:0] Qcoeff[39] = 56;
    reg [7:0] Qcoeff[40] = 49;
    reg [7:0] Qcoeff[41] = 3A;
    reg [7:0] Qcoeff[42] = 2B;
    reg [7:0] Qcoeff[43] = 1D;
    reg [7:0] Qcoeff[44] = 10;
    reg [7:0] Qcoeff[45] = 06;
    reg [7:0] Qcoeff[46] = FE;
    reg [7:0] Qcoeff[47] = F8;
    reg [7:0] Qcoeff[48] = F5;
    reg [7:0] Qcoeff[49] = F4;
    reg [7:0] Qcoeff[50] = F4;
    reg [7:0] Qcoeff[51] = F6;
    reg [7:0] Qcoeff[52] = F9;
    reg [7:0] Qcoeff[53] = FB;
    reg [7:0] Qcoeff[54] = FE;
    reg [7:0] Qcoeff[55] = 01;
    reg [7:0] Qcoeff[56] = 02;
    reg [7:0] Qcoeff[57] = 03;
    reg [7:0] Qcoeff[58] = 03;
    reg [7:0] Qcoeff[59] = 03;
    reg [7:0] Qcoeff[60] = 02;
    reg [7:0] Qcoeff[61] = 00;
    reg [7:0] Qcoeff[62] = FF;
    reg [7:0] Qcoeff[63] = FE;
    reg [7:0] Qcoeff[64] = FE;
    reg [7:0] Qcoeff[65] = FD;
    reg [7:0] Qcoeff[66] = FE;
    reg [7:0] Qcoeff[67] = FE;
    reg [7:0] Qcoeff[68] = FF;
    reg [7:0] Qcoeff[69] = 00;
    reg [7:0] Qcoeff[70] = 00;


    // Transmit Datastream with header
    reg [779:768] datastream = B38;
    reg [767:752] datastream = D196;
    reg [751:736] datastream = 7592;
    reg [735:720] datastream = FAE7;
    reg [719:704] datastream = 8104;
    reg [703:688] datastream = 35D3;
    reg [687:672] datastream = 6897;
    reg [671:656] datastream = 9BF2;
    reg [655:640] datastream = A590;
    reg [639:624] datastream = 451B;
    reg [623:608] datastream = E113;
    reg [607:592] datastream = 15AC;
    reg [591:576] datastream = CB73;
    reg [575:560] datastream = DEBF;
    reg [559:544] datastream = 0193;
    reg [543:528] datastream = 6465;
    reg [527:512] datastream = 02F3;
    reg [511:496] datastream = 9786;
    reg [495:480] datastream = 4A79;
    reg [479:464] datastream = 6B6F;
    reg [463:448] datastream = 2E55;
    reg [447:432] datastream = CDA6;
    reg [431:416] datastream = 8028;
    reg [415:400] datastream = 5FE6;
    reg [399:384] datastream = 80E7;
    reg [383:368] datastream = FE45;
    reg [367:352] datastream = 8CF6;
    reg [351:336] datastream = C49A;
    reg [335:320] datastream = 4E25;
    reg [319:304] datastream = F8C8;
    reg [303:288] datastream = 0985;
    reg [287:272] datastream = FC5F;
    reg [271:256] datastream = 23B5;
    reg [255:240] datastream = 94F7;
    reg [239:224] datastream = B931;
    reg [223:208] datastream = E1FA;
    reg [207:192] datastream = 6604;
    reg [191:176] datastream = CB9A;
    reg [175:160] datastream = EA5C;
    reg [159:144] datastream = 2DE4;
    reg [143:128] datastream = F7BA;
    reg [127:112] datastream = 962F;
    reg [111:96] datastream = 329D;
    reg [95:80] datastream = 7727;
    reg [79:64] datastream = 9533;
    reg [63:48] datastream = 2149;
    reg [47:32] datastream = 386A;
    reg [31:16] datastream = E179;
    reg [15:0] datastream = AA26;


    // I Channel 10b Expected output
    reg [9:0] I_filtered_10b[1733] = 000;
    reg [9:0] I_filtered_10b[1732] = 000;
    reg [9:0] I_filtered_10b[1731] = 000;
    reg [9:0] I_filtered_10b[1730] = 000;
    reg [9:0] I_filtered_10b[1729] = 000;
    reg [9:0] I_filtered_10b[1728] = 000;
    reg [9:0] I_filtered_10b[1727] = 000;
    reg [9:0] I_filtered_10b[1726] = 000;
    reg [9:0] I_filtered_10b[1725] = 000;
    reg [9:0] I_filtered_10b[1724] = 000;
    reg [9:0] I_filtered_10b[1723] = 000;
    reg [9:0] I_filtered_10b[1722] = 000;
    reg [9:0] I_filtered_10b[1721] = 000;
    reg [9:0] I_filtered_10b[1720] = 000;
    reg [9:0] I_filtered_10b[1719] = 000;
    reg [9:0] I_filtered_10b[1718] = 000;
    reg [9:0] I_filtered_10b[1717] = 000;
    reg [9:0] I_filtered_10b[1716] = 001;
    reg [9:0] I_filtered_10b[1715] = 000;
    reg [9:0] I_filtered_10b[1714] = 000;
    reg [9:0] I_filtered_10b[1713] = 000;
    reg [9:0] I_filtered_10b[1712] = 000;
    reg [9:0] I_filtered_10b[1711] = 000;
    reg [9:0] I_filtered_10b[1710] = 3FF;
    reg [9:0] I_filtered_10b[1709] = 3FF;
    reg [9:0] I_filtered_10b[1708] = 3FF;
    reg [9:0] I_filtered_10b[1707] = 000;
    reg [9:0] I_filtered_10b[1706] = 001;
    reg [9:0] I_filtered_10b[1705] = 004;
    reg [9:0] I_filtered_10b[1704] = 005;
    reg [9:0] I_filtered_10b[1703] = 007;
    reg [9:0] I_filtered_10b[1702] = 006;
    reg [9:0] I_filtered_10b[1701] = 007;
    reg [9:0] I_filtered_10b[1700] = 005;
    reg [9:0] I_filtered_10b[1699] = 003;
    reg [9:0] I_filtered_10b[1698] = 3FF;
    reg [9:0] I_filtered_10b[1697] = 3FB;
    reg [9:0] I_filtered_10b[1696] = 3F9;
    reg [9:0] I_filtered_10b[1695] = 3F6;
    reg [9:0] I_filtered_10b[1694] = 3F5;
    reg [9:0] I_filtered_10b[1693] = 3F3;
    reg [9:0] I_filtered_10b[1692] = 3F5;
    reg [9:0] I_filtered_10b[1691] = 3F6;
    reg [9:0] I_filtered_10b[1690] = 3F8;
    reg [9:0] I_filtered_10b[1689] = 3FA;
    reg [9:0] I_filtered_10b[1688] = 3FB;
    reg [9:0] I_filtered_10b[1687] = 3F8;
    reg [9:0] I_filtered_10b[1686] = 3F5;
    reg [9:0] I_filtered_10b[1685] = 3EF;
    reg [9:0] I_filtered_10b[1684] = 3E4;
    reg [9:0] I_filtered_10b[1683] = 3D6;
    reg [9:0] I_filtered_10b[1682] = 3C6;
    reg [9:0] I_filtered_10b[1681] = 3B2;
    reg [9:0] I_filtered_10b[1680] = 39C;
    reg [9:0] I_filtered_10b[1679] = 386;
    reg [9:0] I_filtered_10b[1678] = 36F;
    reg [9:0] I_filtered_10b[1677] = 35A;
    reg [9:0] I_filtered_10b[1676] = 348;
    reg [9:0] I_filtered_10b[1675] = 33B;
    reg [9:0] I_filtered_10b[1674] = 332;
    reg [9:0] I_filtered_10b[1673] = 32E;
    reg [9:0] I_filtered_10b[1672] = 32F;
    reg [9:0] I_filtered_10b[1671] = 334;
    reg [9:0] I_filtered_10b[1670] = 33E;
    reg [9:0] I_filtered_10b[1669] = 34C;
    reg [9:0] I_filtered_10b[1668] = 35B;
    reg [9:0] I_filtered_10b[1667] = 36C;
    reg [9:0] I_filtered_10b[1666] = 37C;
    reg [9:0] I_filtered_10b[1665] = 38C;
    reg [9:0] I_filtered_10b[1664] = 399;
    reg [9:0] I_filtered_10b[1663] = 3A4;
    reg [9:0] I_filtered_10b[1662] = 3AC;
    reg [9:0] I_filtered_10b[1661] = 3B5;
    reg [9:0] I_filtered_10b[1660] = 3B9;
    reg [9:0] I_filtered_10b[1659] = 3BC;
    reg [9:0] I_filtered_10b[1658] = 3BF;
    reg [9:0] I_filtered_10b[1657] = 3C1;
    reg [9:0] I_filtered_10b[1656] = 3C3;
    reg [9:0] I_filtered_10b[1655] = 3C5;
    reg [9:0] I_filtered_10b[1654] = 3C7;
    reg [9:0] I_filtered_10b[1653] = 3C8;
    reg [9:0] I_filtered_10b[1652] = 3CD;
    reg [9:0] I_filtered_10b[1651] = 3D0;
    reg [9:0] I_filtered_10b[1650] = 3D5;
    reg [9:0] I_filtered_10b[1649] = 3D9;
    reg [9:0] I_filtered_10b[1648] = 3E0;
    reg [9:0] I_filtered_10b[1647] = 3E6;
    reg [9:0] I_filtered_10b[1646] = 3ED;
    reg [9:0] I_filtered_10b[1645] = 3F3;
    reg [9:0] I_filtered_10b[1644] = 3F6;
    reg [9:0] I_filtered_10b[1643] = 3FC;
    reg [9:0] I_filtered_10b[1642] = 3FE;
    reg [9:0] I_filtered_10b[1641] = 002;
    reg [9:0] I_filtered_10b[1640] = 003;
    reg [9:0] I_filtered_10b[1639] = 005;
    reg [9:0] I_filtered_10b[1638] = 008;
    reg [9:0] I_filtered_10b[1637] = 00A;
    reg [9:0] I_filtered_10b[1636] = 00C;
    reg [9:0] I_filtered_10b[1635] = 010;
    reg [9:0] I_filtered_10b[1634] = 014;
    reg [9:0] I_filtered_10b[1633] = 017;
    reg [9:0] I_filtered_10b[1632] = 01F;
    reg [9:0] I_filtered_10b[1631] = 027;
    reg [9:0] I_filtered_10b[1630] = 032;
    reg [9:0] I_filtered_10b[1629] = 03E;
    reg [9:0] I_filtered_10b[1628] = 04E;
    reg [9:0] I_filtered_10b[1627] = 05D;
    reg [9:0] I_filtered_10b[1626] = 06E;
    reg [9:0] I_filtered_10b[1625] = 07E;
    reg [9:0] I_filtered_10b[1624] = 08C;
    reg [9:0] I_filtered_10b[1623] = 097;
    reg [9:0] I_filtered_10b[1622] = 09D;
    reg [9:0] I_filtered_10b[1621] = 09F;
    reg [9:0] I_filtered_10b[1620] = 09B;
    reg [9:0] I_filtered_10b[1619] = 092;
    reg [9:0] I_filtered_10b[1618] = 083;
    reg [9:0] I_filtered_10b[1617] = 071;
    reg [9:0] I_filtered_10b[1616] = 05C;
    reg [9:0] I_filtered_10b[1615] = 043;
    reg [9:0] I_filtered_10b[1614] = 02C;
    reg [9:0] I_filtered_10b[1613] = 015;
    reg [9:0] I_filtered_10b[1612] = 000;
    reg [9:0] I_filtered_10b[1611] = 3F1;
    reg [9:0] I_filtered_10b[1610] = 3E3;
    reg [9:0] I_filtered_10b[1609] = 3D9;
    reg [9:0] I_filtered_10b[1608] = 3D4;
    reg [9:0] I_filtered_10b[1607] = 3D3;
    reg [9:0] I_filtered_10b[1606] = 3D3;
    reg [9:0] I_filtered_10b[1605] = 3D6;
    reg [9:0] I_filtered_10b[1604] = 3DA;
    reg [9:0] I_filtered_10b[1603] = 3DE;
    reg [9:0] I_filtered_10b[1602] = 3E1;
    reg [9:0] I_filtered_10b[1601] = 3E3;
    reg [9:0] I_filtered_10b[1600] = 3E4;
    reg [9:0] I_filtered_10b[1599] = 3E3;
    reg [9:0] I_filtered_10b[1598] = 3E3;
    reg [9:0] I_filtered_10b[1597] = 3E2;
    reg [9:0] I_filtered_10b[1596] = 3E2;
    reg [9:0] I_filtered_10b[1595] = 3E0;
    reg [9:0] I_filtered_10b[1594] = 3E2;
    reg [9:0] I_filtered_10b[1593] = 3E5;
    reg [9:0] I_filtered_10b[1592] = 3E9;
    reg [9:0] I_filtered_10b[1591] = 3ED;
    reg [9:0] I_filtered_10b[1590] = 3F4;
    reg [9:0] I_filtered_10b[1589] = 3FC;
    reg [9:0] I_filtered_10b[1588] = 002;
    reg [9:0] I_filtered_10b[1587] = 009;
    reg [9:0] I_filtered_10b[1586] = 00F;
    reg [9:0] I_filtered_10b[1585] = 012;
    reg [9:0] I_filtered_10b[1584] = 015;
    reg [9:0] I_filtered_10b[1583] = 018;
    reg [9:0] I_filtered_10b[1582] = 01A;
    reg [9:0] I_filtered_10b[1581] = 01A;
    reg [9:0] I_filtered_10b[1580] = 01E;
    reg [9:0] I_filtered_10b[1579] = 021;
    reg [9:0] I_filtered_10b[1578] = 026;
    reg [9:0] I_filtered_10b[1577] = 02C;
    reg [9:0] I_filtered_10b[1576] = 035;
    reg [9:0] I_filtered_10b[1575] = 040;
    reg [9:0] I_filtered_10b[1574] = 04A;
    reg [9:0] I_filtered_10b[1573] = 055;
    reg [9:0] I_filtered_10b[1572] = 05D;
    reg [9:0] I_filtered_10b[1571] = 064;
    reg [9:0] I_filtered_10b[1570] = 066;
    reg [9:0] I_filtered_10b[1569] = 065;
    reg [9:0] I_filtered_10b[1568] = 05F;
    reg [9:0] I_filtered_10b[1567] = 054;
    reg [9:0] I_filtered_10b[1566] = 046;
    reg [9:0] I_filtered_10b[1565] = 035;
    reg [9:0] I_filtered_10b[1564] = 021;
    reg [9:0] I_filtered_10b[1563] = 00A;
    reg [9:0] I_filtered_10b[1562] = 3F6;
    reg [9:0] I_filtered_10b[1561] = 3E1;
    reg [9:0] I_filtered_10b[1560] = 3CE;
    reg [9:0] I_filtered_10b[1559] = 3C1;
    reg [9:0] I_filtered_10b[1558] = 3B5;
    reg [9:0] I_filtered_10b[1557] = 3AC;
    reg [9:0] I_filtered_10b[1556] = 3A7;
    reg [9:0] I_filtered_10b[1555] = 3A5;
    reg [9:0] I_filtered_10b[1554] = 3A1;
    reg [9:0] I_filtered_10b[1553] = 39F;
    reg [9:0] I_filtered_10b[1552] = 39D;
    reg [9:0] I_filtered_10b[1551] = 399;
    reg [9:0] I_filtered_10b[1550] = 393;
    reg [9:0] I_filtered_10b[1549] = 38C;
    reg [9:0] I_filtered_10b[1548] = 381;
    reg [9:0] I_filtered_10b[1547] = 378;
    reg [9:0] I_filtered_10b[1546] = 36D;
    reg [9:0] I_filtered_10b[1545] = 366;
    reg [9:0] I_filtered_10b[1544] = 363;
    reg [9:0] I_filtered_10b[1543] = 361;
    reg [9:0] I_filtered_10b[1542] = 366;
    reg [9:0] I_filtered_10b[1541] = 371;
    reg [9:0] I_filtered_10b[1540] = 383;
    reg [9:0] I_filtered_10b[1539] = 399;
    reg [9:0] I_filtered_10b[1538] = 3B5;
    reg [9:0] I_filtered_10b[1537] = 3D5;
    reg [9:0] I_filtered_10b[1536] = 3F5;
    reg [9:0] I_filtered_10b[1535] = 016;
    reg [9:0] I_filtered_10b[1534] = 033;
    reg [9:0] I_filtered_10b[1533] = 04B;
    reg [9:0] I_filtered_10b[1532] = 05E;
    reg [9:0] I_filtered_10b[1531] = 06B;
    reg [9:0] I_filtered_10b[1530] = 071;
    reg [9:0] I_filtered_10b[1529] = 06F;
    reg [9:0] I_filtered_10b[1528] = 069;
    reg [9:0] I_filtered_10b[1527] = 05D;
    reg [9:0] I_filtered_10b[1526] = 04D;
    reg [9:0] I_filtered_10b[1525] = 03B;
    reg [9:0] I_filtered_10b[1524] = 026;
    reg [9:0] I_filtered_10b[1523] = 013;
    reg [9:0] I_filtered_10b[1522] = 003;
    reg [9:0] I_filtered_10b[1521] = 3F6;
    reg [9:0] I_filtered_10b[1520] = 3ED;
    reg [9:0] I_filtered_10b[1519] = 3E5;
    reg [9:0] I_filtered_10b[1518] = 3E1;
    reg [9:0] I_filtered_10b[1517] = 3E0;
    reg [9:0] I_filtered_10b[1516] = 3E1;
    reg [9:0] I_filtered_10b[1515] = 3DF;
    reg [9:0] I_filtered_10b[1514] = 3DC;
    reg [9:0] I_filtered_10b[1513] = 3DB;
    reg [9:0] I_filtered_10b[1512] = 3D4;
    reg [9:0] I_filtered_10b[1511] = 3CD;
    reg [9:0] I_filtered_10b[1510] = 3C3;
    reg [9:0] I_filtered_10b[1509] = 3B8;
    reg [9:0] I_filtered_10b[1508] = 3AE;
    reg [9:0] I_filtered_10b[1507] = 3A5;
    reg [9:0] I_filtered_10b[1506] = 39E;
    reg [9:0] I_filtered_10b[1505] = 39C;
    reg [9:0] I_filtered_10b[1504] = 39B;
    reg [9:0] I_filtered_10b[1503] = 3A0;
    reg [9:0] I_filtered_10b[1502] = 3A9;
    reg [9:0] I_filtered_10b[1501] = 3B7;
    reg [9:0] I_filtered_10b[1500] = 3C8;
    reg [9:0] I_filtered_10b[1499] = 3DD;
    reg [9:0] I_filtered_10b[1498] = 3F5;
    reg [9:0] I_filtered_10b[1497] = 00B;
    reg [9:0] I_filtered_10b[1496] = 022;
    reg [9:0] I_filtered_10b[1495] = 036;
    reg [9:0] I_filtered_10b[1494] = 045;
    reg [9:0] I_filtered_10b[1493] = 052;
    reg [9:0] I_filtered_10b[1492] = 05B;
    reg [9:0] I_filtered_10b[1491] = 05F;
    reg [9:0] I_filtered_10b[1490] = 05F;
    reg [9:0] I_filtered_10b[1489] = 060;
    reg [9:0] I_filtered_10b[1488] = 05D;
    reg [9:0] I_filtered_10b[1487] = 05A;
    reg [9:0] I_filtered_10b[1486] = 057;
    reg [9:0] I_filtered_10b[1485] = 054;
    reg [9:0] I_filtered_10b[1484] = 052;
    reg [9:0] I_filtered_10b[1483] = 054;
    reg [9:0] I_filtered_10b[1482] = 055;
    reg [9:0] I_filtered_10b[1481] = 05A;
    reg [9:0] I_filtered_10b[1480] = 05D;
    reg [9:0] I_filtered_10b[1479] = 05E;
    reg [9:0] I_filtered_10b[1478] = 05F;
    reg [9:0] I_filtered_10b[1477] = 05E;
    reg [9:0] I_filtered_10b[1476] = 056;
    reg [9:0] I_filtered_10b[1475] = 049;
    reg [9:0] I_filtered_10b[1474] = 03A;
    reg [9:0] I_filtered_10b[1473] = 025;
    reg [9:0] I_filtered_10b[1472] = 00C;
    reg [9:0] I_filtered_10b[1471] = 3F1;
    reg [9:0] I_filtered_10b[1470] = 3D4;
    reg [9:0] I_filtered_10b[1469] = 3BA;
    reg [9:0] I_filtered_10b[1468] = 3A6;
    reg [9:0] I_filtered_10b[1467] = 395;
    reg [9:0] I_filtered_10b[1466] = 38C;
    reg [9:0] I_filtered_10b[1465] = 389;
    reg [9:0] I_filtered_10b[1464] = 38F;
    reg [9:0] I_filtered_10b[1463] = 39D;
    reg [9:0] I_filtered_10b[1462] = 3B1;
    reg [9:0] I_filtered_10b[1461] = 3CA;
    reg [9:0] I_filtered_10b[1460] = 3E9;
    reg [9:0] I_filtered_10b[1459] = 00A;
    reg [9:0] I_filtered_10b[1458] = 02A;
    reg [9:0] I_filtered_10b[1457] = 049;
    reg [9:0] I_filtered_10b[1456] = 063;
    reg [9:0] I_filtered_10b[1455] = 078;
    reg [9:0] I_filtered_10b[1454] = 089;
    reg [9:0] I_filtered_10b[1453] = 094;
    reg [9:0] I_filtered_10b[1452] = 099;
    reg [9:0] I_filtered_10b[1451] = 099;
    reg [9:0] I_filtered_10b[1450] = 09A;
    reg [9:0] I_filtered_10b[1449] = 097;
    reg [9:0] I_filtered_10b[1448] = 091;
    reg [9:0] I_filtered_10b[1447] = 08F;
    reg [9:0] I_filtered_10b[1446] = 08C;
    reg [9:0] I_filtered_10b[1445] = 08C;
    reg [9:0] I_filtered_10b[1444] = 08E;
    reg [9:0] I_filtered_10b[1443] = 090;
    reg [9:0] I_filtered_10b[1442] = 093;
    reg [9:0] I_filtered_10b[1441] = 095;
    reg [9:0] I_filtered_10b[1440] = 093;
    reg [9:0] I_filtered_10b[1439] = 093;
    reg [9:0] I_filtered_10b[1438] = 08D;
    reg [9:0] I_filtered_10b[1437] = 084;
    reg [9:0] I_filtered_10b[1436] = 078;
    reg [9:0] I_filtered_10b[1435] = 069;
    reg [9:0] I_filtered_10b[1434] = 057;
    reg [9:0] I_filtered_10b[1433] = 041;
    reg [9:0] I_filtered_10b[1432] = 02D;
    reg [9:0] I_filtered_10b[1431] = 017;
    reg [9:0] I_filtered_10b[1430] = 004;
    reg [9:0] I_filtered_10b[1429] = 3F7;
    reg [9:0] I_filtered_10b[1428] = 3EB;
    reg [9:0] I_filtered_10b[1427] = 3E1;
    reg [9:0] I_filtered_10b[1426] = 3DA;
    reg [9:0] I_filtered_10b[1425] = 3D9;
    reg [9:0] I_filtered_10b[1424] = 3D5;
    reg [9:0] I_filtered_10b[1423] = 3D3;
    reg [9:0] I_filtered_10b[1422] = 3D1;
    reg [9:0] I_filtered_10b[1421] = 3CE;
    reg [9:0] I_filtered_10b[1420] = 3C8;
    reg [9:0] I_filtered_10b[1419] = 3C0;
    reg [9:0] I_filtered_10b[1418] = 3B6;
    reg [9:0] I_filtered_10b[1417] = 3AB;
    reg [9:0] I_filtered_10b[1416] = 3A1;
    reg [9:0] I_filtered_10b[1415] = 399;
    reg [9:0] I_filtered_10b[1414] = 396;
    reg [9:0] I_filtered_10b[1413] = 395;
    reg [9:0] I_filtered_10b[1412] = 39B;
    reg [9:0] I_filtered_10b[1411] = 3A7;
    reg [9:0] I_filtered_10b[1410] = 3BA;
    reg [9:0] I_filtered_10b[1409] = 3CF;
    reg [9:0] I_filtered_10b[1408] = 3EC;
    reg [9:0] I_filtered_10b[1407] = 00C;
    reg [9:0] I_filtered_10b[1406] = 02B;
    reg [9:0] I_filtered_10b[1405] = 04B;
    reg [9:0] I_filtered_10b[1404] = 067;
    reg [9:0] I_filtered_10b[1403] = 07C;
    reg [9:0] I_filtered_10b[1402] = 08E;
    reg [9:0] I_filtered_10b[1401] = 09A;
    reg [9:0] I_filtered_10b[1400] = 09F;
    reg [9:0] I_filtered_10b[1399] = 09D;
    reg [9:0] I_filtered_10b[1398] = 09A;
    reg [9:0] I_filtered_10b[1397] = 092;
    reg [9:0] I_filtered_10b[1396] = 088;
    reg [9:0] I_filtered_10b[1395] = 07F;
    reg [9:0] I_filtered_10b[1394] = 073;
    reg [9:0] I_filtered_10b[1393] = 06A;
    reg [9:0] I_filtered_10b[1392] = 066;
    reg [9:0] I_filtered_10b[1391] = 061;
    reg [9:0] I_filtered_10b[1390] = 062;
    reg [9:0] I_filtered_10b[1389] = 061;
    reg [9:0] I_filtered_10b[1388] = 05F;
    reg [9:0] I_filtered_10b[1387] = 05F;
    reg [9:0] I_filtered_10b[1386] = 05D;
    reg [9:0] I_filtered_10b[1385] = 052;
    reg [9:0] I_filtered_10b[1384] = 042;
    reg [9:0] I_filtered_10b[1383] = 02F;
    reg [9:0] I_filtered_10b[1382] = 013;
    reg [9:0] I_filtered_10b[1381] = 3F6;
    reg [9:0] I_filtered_10b[1380] = 3D4;
    reg [9:0] I_filtered_10b[1379] = 3AE;
    reg [9:0] I_filtered_10b[1378] = 38E;
    reg [9:0] I_filtered_10b[1377] = 36F;
    reg [9:0] I_filtered_10b[1376] = 358;
    reg [9:0] I_filtered_10b[1375] = 34A;
    reg [9:0] I_filtered_10b[1374] = 343;
    reg [9:0] I_filtered_10b[1373] = 348;
    reg [9:0] I_filtered_10b[1372] = 359;
    reg [9:0] I_filtered_10b[1371] = 377;
    reg [9:0] I_filtered_10b[1370] = 39C;
    reg [9:0] I_filtered_10b[1369] = 3CB;
    reg [9:0] I_filtered_10b[1368] = 3FE;
    reg [9:0] I_filtered_10b[1367] = 031;
    reg [9:0] I_filtered_10b[1366] = 067;
    reg [9:0] I_filtered_10b[1365] = 094;
    reg [9:0] I_filtered_10b[1364] = 0BD;
    reg [9:0] I_filtered_10b[1363] = 0DB;
    reg [9:0] I_filtered_10b[1362] = 0EF;
    reg [9:0] I_filtered_10b[1361] = 0F6;
    reg [9:0] I_filtered_10b[1360] = 0F4;
    reg [9:0] I_filtered_10b[1359] = 0E6;
    reg [9:0] I_filtered_10b[1358] = 0CB;
    reg [9:0] I_filtered_10b[1357] = 0A7;
    reg [9:0] I_filtered_10b[1356] = 07E;
    reg [9:0] I_filtered_10b[1355] = 04F;
    reg [9:0] I_filtered_10b[1354] = 020;
    reg [9:0] I_filtered_10b[1353] = 3F2;
    reg [9:0] I_filtered_10b[1352] = 3C8;
    reg [9:0] I_filtered_10b[1351] = 3A5;
    reg [9:0] I_filtered_10b[1350] = 38A;
    reg [9:0] I_filtered_10b[1349] = 37A;
    reg [9:0] I_filtered_10b[1348] = 377;
    reg [9:0] I_filtered_10b[1347] = 37C;
    reg [9:0] I_filtered_10b[1346] = 38D;
    reg [9:0] I_filtered_10b[1345] = 3A8;
    reg [9:0] I_filtered_10b[1344] = 3CB;
    reg [9:0] I_filtered_10b[1343] = 3F4;
    reg [9:0] I_filtered_10b[1342] = 021;
    reg [9:0] I_filtered_10b[1341] = 04E;
    reg [9:0] I_filtered_10b[1340] = 07A;
    reg [9:0] I_filtered_10b[1339] = 0A2;
    reg [9:0] I_filtered_10b[1338] = 0C4;
    reg [9:0] I_filtered_10b[1337] = 0DE;
    reg [9:0] I_filtered_10b[1336] = 0ED;
    reg [9:0] I_filtered_10b[1335] = 0F0;
    reg [9:0] I_filtered_10b[1334] = 0EC;
    reg [9:0] I_filtered_10b[1333] = 0DC;
    reg [9:0] I_filtered_10b[1332] = 0C2;
    reg [9:0] I_filtered_10b[1331] = 09F;
    reg [9:0] I_filtered_10b[1330] = 078;
    reg [9:0] I_filtered_10b[1329] = 04B;
    reg [9:0] I_filtered_10b[1328] = 01E;
    reg [9:0] I_filtered_10b[1327] = 3F3;
    reg [9:0] I_filtered_10b[1326] = 3CB;
    reg [9:0] I_filtered_10b[1325] = 3AA;
    reg [9:0] I_filtered_10b[1324] = 390;
    reg [9:0] I_filtered_10b[1323] = 381;
    reg [9:0] I_filtered_10b[1322] = 37D;
    reg [9:0] I_filtered_10b[1321] = 382;
    reg [9:0] I_filtered_10b[1320] = 390;
    reg [9:0] I_filtered_10b[1319] = 3A6;
    reg [9:0] I_filtered_10b[1318] = 3C4;
    reg [9:0] I_filtered_10b[1317] = 3E5;
    reg [9:0] I_filtered_10b[1316] = 00B;
    reg [9:0] I_filtered_10b[1315] = 02F;
    reg [9:0] I_filtered_10b[1314] = 051;
    reg [9:0] I_filtered_10b[1313] = 070;
    reg [9:0] I_filtered_10b[1312] = 087;
    reg [9:0] I_filtered_10b[1311] = 09A;
    reg [9:0] I_filtered_10b[1310] = 0A4;
    reg [9:0] I_filtered_10b[1309] = 0A5;
    reg [9:0] I_filtered_10b[1308] = 0A0;
    reg [9:0] I_filtered_10b[1307] = 098;
    reg [9:0] I_filtered_10b[1306] = 08C;
    reg [9:0] I_filtered_10b[1305] = 07B;
    reg [9:0] I_filtered_10b[1304] = 06C;
    reg [9:0] I_filtered_10b[1303] = 05A;
    reg [9:0] I_filtered_10b[1302] = 04D;
    reg [9:0] I_filtered_10b[1301] = 041;
    reg [9:0] I_filtered_10b[1300] = 036;
    reg [9:0] I_filtered_10b[1299] = 02C;
    reg [9:0] I_filtered_10b[1298] = 025;
    reg [9:0] I_filtered_10b[1297] = 01D;
    reg [9:0] I_filtered_10b[1296] = 01A;
    reg [9:0] I_filtered_10b[1295] = 014;
    reg [9:0] I_filtered_10b[1294] = 00D;
    reg [9:0] I_filtered_10b[1293] = 006;
    reg [9:0] I_filtered_10b[1292] = 3FF;
    reg [9:0] I_filtered_10b[1291] = 3F5;
    reg [9:0] I_filtered_10b[1290] = 3EC;
    reg [9:0] I_filtered_10b[1289] = 3E4;
    reg [9:0] I_filtered_10b[1288] = 3D8;
    reg [9:0] I_filtered_10b[1287] = 3D0;
    reg [9:0] I_filtered_10b[1286] = 3C5;
    reg [9:0] I_filtered_10b[1285] = 3BE;
    reg [9:0] I_filtered_10b[1284] = 3B5;
    reg [9:0] I_filtered_10b[1283] = 3AD;
    reg [9:0] I_filtered_10b[1282] = 3A6;
    reg [9:0] I_filtered_10b[1281] = 39E;
    reg [9:0] I_filtered_10b[1280] = 39B;
    reg [9:0] I_filtered_10b[1279] = 397;
    reg [9:0] I_filtered_10b[1278] = 394;
    reg [9:0] I_filtered_10b[1277] = 390;
    reg [9:0] I_filtered_10b[1276] = 38F;
    reg [9:0] I_filtered_10b[1275] = 38D;
    reg [9:0] I_filtered_10b[1274] = 38A;
    reg [9:0] I_filtered_10b[1273] = 387;
    reg [9:0] I_filtered_10b[1272] = 385;
    reg [9:0] I_filtered_10b[1271] = 382;
    reg [9:0] I_filtered_10b[1270] = 37F;
    reg [9:0] I_filtered_10b[1269] = 37D;
    reg [9:0] I_filtered_10b[1268] = 377;
    reg [9:0] I_filtered_10b[1267] = 373;
    reg [9:0] I_filtered_10b[1266] = 36D;
    reg [9:0] I_filtered_10b[1265] = 366;
    reg [9:0] I_filtered_10b[1264] = 35D;
    reg [9:0] I_filtered_10b[1263] = 354;
    reg [9:0] I_filtered_10b[1262] = 34B;
    reg [9:0] I_filtered_10b[1261] = 342;
    reg [9:0] I_filtered_10b[1260] = 33A;
    reg [9:0] I_filtered_10b[1259] = 334;
    reg [9:0] I_filtered_10b[1258] = 333;
    reg [9:0] I_filtered_10b[1257] = 334;
    reg [9:0] I_filtered_10b[1256] = 338;
    reg [9:0] I_filtered_10b[1255] = 341;
    reg [9:0] I_filtered_10b[1254] = 34E;
    reg [9:0] I_filtered_10b[1253] = 35F;
    reg [9:0] I_filtered_10b[1252] = 372;
    reg [9:0] I_filtered_10b[1251] = 388;
    reg [9:0] I_filtered_10b[1250] = 39C;
    reg [9:0] I_filtered_10b[1249] = 3B2;
    reg [9:0] I_filtered_10b[1248] = 3C6;
    reg [9:0] I_filtered_10b[1247] = 3D7;
    reg [9:0] I_filtered_10b[1246] = 3E5;
    reg [9:0] I_filtered_10b[1245] = 3F1;
    reg [9:0] I_filtered_10b[1244] = 3F8;
    reg [9:0] I_filtered_10b[1243] = 3FC;
    reg [9:0] I_filtered_10b[1242] = 3FD;
    reg [9:0] I_filtered_10b[1241] = 3FA;
    reg [9:0] I_filtered_10b[1240] = 3F6;
    reg [9:0] I_filtered_10b[1239] = 3F0;
    reg [9:0] I_filtered_10b[1238] = 3E9;
    reg [9:0] I_filtered_10b[1237] = 3E0;
    reg [9:0] I_filtered_10b[1236] = 3DC;
    reg [9:0] I_filtered_10b[1235] = 3D7;
    reg [9:0] I_filtered_10b[1234] = 3D8;
    reg [9:0] I_filtered_10b[1233] = 3D7;
    reg [9:0] I_filtered_10b[1232] = 3DB;
    reg [9:0] I_filtered_10b[1231] = 3E0;
    reg [9:0] I_filtered_10b[1230] = 3E7;
    reg [9:0] I_filtered_10b[1229] = 3EE;
    reg [9:0] I_filtered_10b[1228] = 3F2;
    reg [9:0] I_filtered_10b[1227] = 3F9;
    reg [9:0] I_filtered_10b[1226] = 3FC;
    reg [9:0] I_filtered_10b[1225] = 000;
    reg [9:0] I_filtered_10b[1224] = 000;
    reg [9:0] I_filtered_10b[1223] = 000;
    reg [9:0] I_filtered_10b[1222] = 001;
    reg [9:0] I_filtered_10b[1221] = 003;
    reg [9:0] I_filtered_10b[1220] = 004;
    reg [9:0] I_filtered_10b[1219] = 009;
    reg [9:0] I_filtered_10b[1218] = 00E;
    reg [9:0] I_filtered_10b[1217] = 015;
    reg [9:0] I_filtered_10b[1216] = 022;
    reg [9:0] I_filtered_10b[1215] = 02E;
    reg [9:0] I_filtered_10b[1214] = 03E;
    reg [9:0] I_filtered_10b[1213] = 050;
    reg [9:0] I_filtered_10b[1212] = 066;
    reg [9:0] I_filtered_10b[1211] = 07A;
    reg [9:0] I_filtered_10b[1210] = 08F;
    reg [9:0] I_filtered_10b[1209] = 0A2;
    reg [9:0] I_filtered_10b[1208] = 0B2;
    reg [9:0] I_filtered_10b[1207] = 0BF;
    reg [9:0] I_filtered_10b[1206] = 0C8;
    reg [9:0] I_filtered_10b[1205] = 0CC;
    reg [9:0] I_filtered_10b[1204] = 0CC;
    reg [9:0] I_filtered_10b[1203] = 0CA;
    reg [9:0] I_filtered_10b[1202] = 0C4;
    reg [9:0] I_filtered_10b[1201] = 0BC;
    reg [9:0] I_filtered_10b[1200] = 0B4;
    reg [9:0] I_filtered_10b[1199] = 0AA;
    reg [9:0] I_filtered_10b[1198] = 0A1;
    reg [9:0] I_filtered_10b[1197] = 09B;
    reg [9:0] I_filtered_10b[1196] = 095;
    reg [9:0] I_filtered_10b[1195] = 094;
    reg [9:0] I_filtered_10b[1194] = 092;
    reg [9:0] I_filtered_10b[1193] = 08E;
    reg [9:0] I_filtered_10b[1192] = 08D;
    reg [9:0] I_filtered_10b[1191] = 08B;
    reg [9:0] I_filtered_10b[1190] = 083;
    reg [9:0] I_filtered_10b[1189] = 078;
    reg [9:0] I_filtered_10b[1188] = 06A;
    reg [9:0] I_filtered_10b[1187] = 057;
    reg [9:0] I_filtered_10b[1186] = 040;
    reg [9:0] I_filtered_10b[1185] = 027;
    reg [9:0] I_filtered_10b[1184] = 00C;
    reg [9:0] I_filtered_10b[1183] = 3F2;
    reg [9:0] I_filtered_10b[1182] = 3DD;
    reg [9:0] I_filtered_10b[1181] = 3CC;
    reg [9:0] I_filtered_10b[1180] = 3C1;
    reg [9:0] I_filtered_10b[1179] = 3BC;
    reg [9:0] I_filtered_10b[1178] = 3C2;
    reg [9:0] I_filtered_10b[1177] = 3CF;
    reg [9:0] I_filtered_10b[1176] = 3E4;
    reg [9:0] I_filtered_10b[1175] = 3FC;
    reg [9:0] I_filtered_10b[1174] = 01C;
    reg [9:0] I_filtered_10b[1173] = 03F;
    reg [9:0] I_filtered_10b[1172] = 060;
    reg [9:0] I_filtered_10b[1171] = 081;
    reg [9:0] I_filtered_10b[1170] = 09C;
    reg [9:0] I_filtered_10b[1169] = 0B2;
    reg [9:0] I_filtered_10b[1168] = 0C4;
    reg [9:0] I_filtered_10b[1167] = 0CF;
    reg [9:0] I_filtered_10b[1166] = 0D2;
    reg [9:0] I_filtered_10b[1165] = 0D2;
    reg [9:0] I_filtered_10b[1164] = 0CF;
    reg [9:0] I_filtered_10b[1163] = 0C8;
    reg [9:0] I_filtered_10b[1162] = 0BD;
    reg [9:0] I_filtered_10b[1161] = 0B5;
    reg [9:0] I_filtered_10b[1160] = 0A9;
    reg [9:0] I_filtered_10b[1159] = 0A0;
    reg [9:0] I_filtered_10b[1158] = 09A;
    reg [9:0] I_filtered_10b[1157] = 092;
    reg [9:0] I_filtered_10b[1156] = 08F;
    reg [9:0] I_filtered_10b[1155] = 08C;
    reg [9:0] I_filtered_10b[1154] = 088;
    reg [9:0] I_filtered_10b[1153] = 087;
    reg [9:0] I_filtered_10b[1152] = 085;
    reg [9:0] I_filtered_10b[1151] = 080;
    reg [9:0] I_filtered_10b[1150] = 079;
    reg [9:0] I_filtered_10b[1149] = 071;
    reg [9:0] I_filtered_10b[1148] = 066;
    reg [9:0] I_filtered_10b[1147] = 058;
    reg [9:0] I_filtered_10b[1146] = 04A;
    reg [9:0] I_filtered_10b[1145] = 039;
    reg [9:0] I_filtered_10b[1144] = 02A;
    reg [9:0] I_filtered_10b[1143] = 01E;
    reg [9:0] I_filtered_10b[1142] = 014;
    reg [9:0] I_filtered_10b[1141] = 00C;
    reg [9:0] I_filtered_10b[1140] = 008;
    reg [9:0] I_filtered_10b[1139] = 009;
    reg [9:0] I_filtered_10b[1138] = 00C;
    reg [9:0] I_filtered_10b[1137] = 013;
    reg [9:0] I_filtered_10b[1136] = 01A;
    reg [9:0] I_filtered_10b[1135] = 025;
    reg [9:0] I_filtered_10b[1134] = 030;
    reg [9:0] I_filtered_10b[1133] = 03B;
    reg [9:0] I_filtered_10b[1132] = 043;
    reg [9:0] I_filtered_10b[1131] = 04A;
    reg [9:0] I_filtered_10b[1130] = 04C;
    reg [9:0] I_filtered_10b[1129] = 04F;
    reg [9:0] I_filtered_10b[1128] = 04F;
    reg [9:0] I_filtered_10b[1127] = 04D;
    reg [9:0] I_filtered_10b[1126] = 04B;
    reg [9:0] I_filtered_10b[1125] = 04D;
    reg [9:0] I_filtered_10b[1124] = 051;
    reg [9:0] I_filtered_10b[1123] = 055;
    reg [9:0] I_filtered_10b[1122] = 05E;
    reg [9:0] I_filtered_10b[1121] = 067;
    reg [9:0] I_filtered_10b[1120] = 074;
    reg [9:0] I_filtered_10b[1119] = 082;
    reg [9:0] I_filtered_10b[1118] = 08E;
    reg [9:0] I_filtered_10b[1117] = 09A;
    reg [9:0] I_filtered_10b[1116] = 0A3;
    reg [9:0] I_filtered_10b[1115] = 0A5;
    reg [9:0] I_filtered_10b[1114] = 0A5;
    reg [9:0] I_filtered_10b[1113] = 09F;
    reg [9:0] I_filtered_10b[1112] = 08F;
    reg [9:0] I_filtered_10b[1111] = 079;
    reg [9:0] I_filtered_10b[1110] = 05D;
    reg [9:0] I_filtered_10b[1109] = 03A;
    reg [9:0] I_filtered_10b[1108] = 011;
    reg [9:0] I_filtered_10b[1107] = 3E8;
    reg [9:0] I_filtered_10b[1106] = 3BD;
    reg [9:0] I_filtered_10b[1105] = 396;
    reg [9:0] I_filtered_10b[1104] = 377;
    reg [9:0] I_filtered_10b[1103] = 35E;
    reg [9:0] I_filtered_10b[1102] = 34F;
    reg [9:0] I_filtered_10b[1101] = 349;
    reg [9:0] I_filtered_10b[1100] = 350;
    reg [9:0] I_filtered_10b[1099] = 35D;
    reg [9:0] I_filtered_10b[1098] = 373;
    reg [9:0] I_filtered_10b[1097] = 38F;
    reg [9:0] I_filtered_10b[1096] = 3AF;
    reg [9:0] I_filtered_10b[1095] = 3D1;
    reg [9:0] I_filtered_10b[1094] = 3F0;
    reg [9:0] I_filtered_10b[1093] = 00D;
    reg [9:0] I_filtered_10b[1092] = 025;
    reg [9:0] I_filtered_10b[1091] = 038;
    reg [9:0] I_filtered_10b[1090] = 047;
    reg [9:0] I_filtered_10b[1089] = 054;
    reg [9:0] I_filtered_10b[1088] = 059;
    reg [9:0] I_filtered_10b[1087] = 05E;
    reg [9:0] I_filtered_10b[1086] = 066;
    reg [9:0] I_filtered_10b[1085] = 06B;
    reg [9:0] I_filtered_10b[1084] = 070;
    reg [9:0] I_filtered_10b[1083] = 07A;
    reg [9:0] I_filtered_10b[1082] = 085;
    reg [9:0] I_filtered_10b[1081] = 090;
    reg [9:0] I_filtered_10b[1080] = 0A0;
    reg [9:0] I_filtered_10b[1079] = 0AC;
    reg [9:0] I_filtered_10b[1078] = 0B8;
    reg [9:0] I_filtered_10b[1077] = 0C2;
    reg [9:0] I_filtered_10b[1076] = 0C8;
    reg [9:0] I_filtered_10b[1075] = 0CC;
    reg [9:0] I_filtered_10b[1074] = 0CB;
    reg [9:0] I_filtered_10b[1073] = 0C7;
    reg [9:0] I_filtered_10b[1072] = 0BD;
    reg [9:0] I_filtered_10b[1071] = 0B2;
    reg [9:0] I_filtered_10b[1070] = 0A4;
    reg [9:0] I_filtered_10b[1069] = 096;
    reg [9:0] I_filtered_10b[1068] = 08A;
    reg [9:0] I_filtered_10b[1067] = 07B;
    reg [9:0] I_filtered_10b[1066] = 071;
    reg [9:0] I_filtered_10b[1065] = 066;
    reg [9:0] I_filtered_10b[1064] = 05F;
    reg [9:0] I_filtered_10b[1063] = 054;
    reg [9:0] I_filtered_10b[1062] = 04D;
    reg [9:0] I_filtered_10b[1061] = 045;
    reg [9:0] I_filtered_10b[1060] = 03C;
    reg [9:0] I_filtered_10b[1059] = 036;
    reg [9:0] I_filtered_10b[1058] = 02E;
    reg [9:0] I_filtered_10b[1057] = 027;
    reg [9:0] I_filtered_10b[1056] = 01E;
    reg [9:0] I_filtered_10b[1055] = 01A;
    reg [9:0] I_filtered_10b[1054] = 011;
    reg [9:0] I_filtered_10b[1053] = 00B;
    reg [9:0] I_filtered_10b[1052] = 004;
    reg [9:0] I_filtered_10b[1051] = 3FE;
    reg [9:0] I_filtered_10b[1050] = 3F5;
    reg [9:0] I_filtered_10b[1049] = 3EC;
    reg [9:0] I_filtered_10b[1048] = 3E4;
    reg [9:0] I_filtered_10b[1047] = 3D6;
    reg [9:0] I_filtered_10b[1046] = 3CB;
    reg [9:0] I_filtered_10b[1045] = 3BB;
    reg [9:0] I_filtered_10b[1044] = 3AB;
    reg [9:0] I_filtered_10b[1043] = 398;
    reg [9:0] I_filtered_10b[1042] = 388;
    reg [9:0] I_filtered_10b[1041] = 373;
    reg [9:0] I_filtered_10b[1040] = 361;
    reg [9:0] I_filtered_10b[1039] = 34E;
    reg [9:0] I_filtered_10b[1038] = 340;
    reg [9:0] I_filtered_10b[1037] = 335;
    reg [9:0] I_filtered_10b[1036] = 32E;
    reg [9:0] I_filtered_10b[1035] = 32B;
    reg [9:0] I_filtered_10b[1034] = 32E;
    reg [9:0] I_filtered_10b[1033] = 338;
    reg [9:0] I_filtered_10b[1032] = 345;
    reg [9:0] I_filtered_10b[1031] = 357;
    reg [9:0] I_filtered_10b[1030] = 368;
    reg [9:0] I_filtered_10b[1029] = 37B;
    reg [9:0] I_filtered_10b[1028] = 390;
    reg [9:0] I_filtered_10b[1027] = 3A1;
    reg [9:0] I_filtered_10b[1026] = 3B1;
    reg [9:0] I_filtered_10b[1025] = 3BD;
    reg [9:0] I_filtered_10b[1024] = 3C7;
    reg [9:0] I_filtered_10b[1023] = 3CB;
    reg [9:0] I_filtered_10b[1022] = 3CD;
    reg [9:0] I_filtered_10b[1021] = 3C7;
    reg [9:0] I_filtered_10b[1020] = 3BB;
    reg [9:0] I_filtered_10b[1019] = 3AD;
    reg [9:0] I_filtered_10b[1018] = 398;
    reg [9:0] I_filtered_10b[1017] = 383;
    reg [9:0] I_filtered_10b[1016] = 369;
    reg [9:0] I_filtered_10b[1015] = 350;
    reg [9:0] I_filtered_10b[1014] = 33A;
    reg [9:0] I_filtered_10b[1013] = 325;
    reg [9:0] I_filtered_10b[1012] = 317;
    reg [9:0] I_filtered_10b[1011] = 313;
    reg [9:0] I_filtered_10b[1010] = 316;
    reg [9:0] I_filtered_10b[1009] = 320;
    reg [9:0] I_filtered_10b[1008] = 337;
    reg [9:0] I_filtered_10b[1007] = 357;
    reg [9:0] I_filtered_10b[1006] = 381;
    reg [9:0] I_filtered_10b[1005] = 3B0;
    reg [9:0] I_filtered_10b[1004] = 3E7;
    reg [9:0] I_filtered_10b[1003] = 01C;
    reg [9:0] I_filtered_10b[1002] = 055;
    reg [9:0] I_filtered_10b[1001] = 088;
    reg [9:0] I_filtered_10b[1000] = 0B6;
    reg [9:0] I_filtered_10b[999] = 0D9;
    reg [9:0] I_filtered_10b[998] = 0F1;
    reg [9:0] I_filtered_10b[997] = 0FC;
    reg [9:0] I_filtered_10b[996] = 0FB;
    reg [9:0] I_filtered_10b[995] = 0EE;
    reg [9:0] I_filtered_10b[994] = 0D2;
    reg [9:0] I_filtered_10b[993] = 0AE;
    reg [9:0] I_filtered_10b[992] = 082;
    reg [9:0] I_filtered_10b[991] = 053;
    reg [9:0] I_filtered_10b[990] = 022;
    reg [9:0] I_filtered_10b[989] = 3F3;
    reg [9:0] I_filtered_10b[988] = 3CB;
    reg [9:0] I_filtered_10b[987] = 3A9;
    reg [9:0] I_filtered_10b[986] = 38F;
    reg [9:0] I_filtered_10b[985] = 380;
    reg [9:0] I_filtered_10b[984] = 37D;
    reg [9:0] I_filtered_10b[983] = 381;
    reg [9:0] I_filtered_10b[982] = 38F;
    reg [9:0] I_filtered_10b[981] = 3A5;
    reg [9:0] I_filtered_10b[980] = 3C4;
    reg [9:0] I_filtered_10b[979] = 3E5;
    reg [9:0] I_filtered_10b[978] = 00C;
    reg [9:0] I_filtered_10b[977] = 032;
    reg [9:0] I_filtered_10b[976] = 056;
    reg [9:0] I_filtered_10b[975] = 078;
    reg [9:0] I_filtered_10b[974] = 092;
    reg [9:0] I_filtered_10b[973] = 0A7;
    reg [9:0] I_filtered_10b[972] = 0B1;
    reg [9:0] I_filtered_10b[971] = 0B1;
    reg [9:0] I_filtered_10b[970] = 0A9;
    reg [9:0] I_filtered_10b[969] = 09A;
    reg [9:0] I_filtered_10b[968] = 085;
    reg [9:0] I_filtered_10b[967] = 069;
    reg [9:0] I_filtered_10b[966] = 04C;
    reg [9:0] I_filtered_10b[965] = 02A;
    reg [9:0] I_filtered_10b[964] = 00D;
    reg [9:0] I_filtered_10b[963] = 3F0;
    reg [9:0] I_filtered_10b[962] = 3D6;
    reg [9:0] I_filtered_10b[961] = 3C0;
    reg [9:0] I_filtered_10b[960] = 3AE;
    reg [9:0] I_filtered_10b[959] = 3A1;
    reg [9:0] I_filtered_10b[958] = 39B;
    reg [9:0] I_filtered_10b[957] = 397;
    reg [9:0] I_filtered_10b[956] = 396;
    reg [9:0] I_filtered_10b[955] = 399;
    reg [9:0] I_filtered_10b[954] = 39F;
    reg [9:0] I_filtered_10b[953] = 3A4;
    reg [9:0] I_filtered_10b[952] = 3A9;
    reg [9:0] I_filtered_10b[951] = 3AF;
    reg [9:0] I_filtered_10b[950] = 3B3;
    reg [9:0] I_filtered_10b[949] = 3B6;
    reg [9:0] I_filtered_10b[948] = 3B9;
    reg [9:0] I_filtered_10b[947] = 3BB;
    reg [9:0] I_filtered_10b[946] = 3BB;
    reg [9:0] I_filtered_10b[945] = 3B9;
    reg [9:0] I_filtered_10b[944] = 3B8;
    reg [9:0] I_filtered_10b[943] = 3B3;
    reg [9:0] I_filtered_10b[942] = 3AE;
    reg [9:0] I_filtered_10b[941] = 3A6;
    reg [9:0] I_filtered_10b[940] = 39E;
    reg [9:0] I_filtered_10b[939] = 395;
    reg [9:0] I_filtered_10b[938] = 38B;
    reg [9:0] I_filtered_10b[937] = 380;
    reg [9:0] I_filtered_10b[936] = 376;
    reg [9:0] I_filtered_10b[935] = 36B;
    reg [9:0] I_filtered_10b[934] = 363;
    reg [9:0] I_filtered_10b[933] = 361;
    reg [9:0] I_filtered_10b[932] = 361;
    reg [9:0] I_filtered_10b[931] = 365;
    reg [9:0] I_filtered_10b[930] = 371;
    reg [9:0] I_filtered_10b[929] = 383;
    reg [9:0] I_filtered_10b[928] = 39A;
    reg [9:0] I_filtered_10b[927] = 3B6;
    reg [9:0] I_filtered_10b[926] = 3D6;
    reg [9:0] I_filtered_10b[925] = 3F7;
    reg [9:0] I_filtered_10b[924] = 01A;
    reg [9:0] I_filtered_10b[923] = 03A;
    reg [9:0] I_filtered_10b[922] = 055;
    reg [9:0] I_filtered_10b[921] = 06A;
    reg [9:0] I_filtered_10b[920] = 078;
    reg [9:0] I_filtered_10b[919] = 07D;
    reg [9:0] I_filtered_10b[918] = 079;
    reg [9:0] I_filtered_10b[917] = 06D;
    reg [9:0] I_filtered_10b[916] = 057;
    reg [9:0] I_filtered_10b[915] = 03D;
    reg [9:0] I_filtered_10b[914] = 01C;
    reg [9:0] I_filtered_10b[913] = 3F9;
    reg [9:0] I_filtered_10b[912] = 3D7;
    reg [9:0] I_filtered_10b[911] = 3B4;
    reg [9:0] I_filtered_10b[910] = 398;
    reg [9:0] I_filtered_10b[909] = 37F;
    reg [9:0] I_filtered_10b[908] = 36C;
    reg [9:0] I_filtered_10b[907] = 35F;
    reg [9:0] I_filtered_10b[906] = 35B;
    reg [9:0] I_filtered_10b[905] = 35B;
    reg [9:0] I_filtered_10b[904] = 361;
    reg [9:0] I_filtered_10b[903] = 36D;
    reg [9:0] I_filtered_10b[902] = 37E;
    reg [9:0] I_filtered_10b[901] = 38F;
    reg [9:0] I_filtered_10b[900] = 3A2;
    reg [9:0] I_filtered_10b[899] = 3B5;
    reg [9:0] I_filtered_10b[898] = 3C8;
    reg [9:0] I_filtered_10b[897] = 3D9;
    reg [9:0] I_filtered_10b[896] = 3E9;
    reg [9:0] I_filtered_10b[895] = 3F4;
    reg [9:0] I_filtered_10b[894] = 3FC;
    reg [9:0] I_filtered_10b[893] = 3FE;
    reg [9:0] I_filtered_10b[892] = 3FF;
    reg [9:0] I_filtered_10b[891] = 3F9;
    reg [9:0] I_filtered_10b[890] = 3EE;
    reg [9:0] I_filtered_10b[889] = 3DF;
    reg [9:0] I_filtered_10b[888] = 3CC;
    reg [9:0] I_filtered_10b[887] = 3B5;
    reg [9:0] I_filtered_10b[886] = 39B;
    reg [9:0] I_filtered_10b[885] = 384;
    reg [9:0] I_filtered_10b[884] = 36D;
    reg [9:0] I_filtered_10b[883] = 35C;
    reg [9:0] I_filtered_10b[882] = 34E;
    reg [9:0] I_filtered_10b[881] = 34B;
    reg [9:0] I_filtered_10b[880] = 34F;
    reg [9:0] I_filtered_10b[879] = 35C;
    reg [9:0] I_filtered_10b[878] = 373;
    reg [9:0] I_filtered_10b[877] = 38F;
    reg [9:0] I_filtered_10b[876] = 3B3;
    reg [9:0] I_filtered_10b[875] = 3DA;
    reg [9:0] I_filtered_10b[874] = 007;
    reg [9:0] I_filtered_10b[873] = 02F;
    reg [9:0] I_filtered_10b[872] = 05A;
    reg [9:0] I_filtered_10b[871] = 07F;
    reg [9:0] I_filtered_10b[870] = 09F;
    reg [9:0] I_filtered_10b[869] = 0B9;
    reg [9:0] I_filtered_10b[868] = 0CD;
    reg [9:0] I_filtered_10b[867] = 0D8;
    reg [9:0] I_filtered_10b[866] = 0DE;
    reg [9:0] I_filtered_10b[865] = 0E1;
    reg [9:0] I_filtered_10b[864] = 0DD;
    reg [9:0] I_filtered_10b[863] = 0D6;
    reg [9:0] I_filtered_10b[862] = 0CF;
    reg [9:0] I_filtered_10b[861] = 0CA;
    reg [9:0] I_filtered_10b[860] = 0C4;
    reg [9:0] I_filtered_10b[859] = 0C0;
    reg [9:0] I_filtered_10b[858] = 0BF;
    reg [9:0] I_filtered_10b[857] = 0BD;
    reg [9:0] I_filtered_10b[856] = 0BC;
    reg [9:0] I_filtered_10b[855] = 0BA;
    reg [9:0] I_filtered_10b[854] = 0BA;
    reg [9:0] I_filtered_10b[853] = 0B6;
    reg [9:0] I_filtered_10b[852] = 0B4;
    reg [9:0] I_filtered_10b[851] = 0B1;
    reg [9:0] I_filtered_10b[850] = 0AF;
    reg [9:0] I_filtered_10b[849] = 0AC;
    reg [9:0] I_filtered_10b[848] = 0A9;
    reg [9:0] I_filtered_10b[847] = 0AA;
    reg [9:0] I_filtered_10b[846] = 0A9;
    reg [9:0] I_filtered_10b[845] = 0AA;
    reg [9:0] I_filtered_10b[844] = 0AC;
    reg [9:0] I_filtered_10b[843] = 0AD;
    reg [9:0] I_filtered_10b[842] = 0A6;
    reg [9:0] I_filtered_10b[841] = 09F;
    reg [9:0] I_filtered_10b[840] = 094;
    reg [9:0] I_filtered_10b[839] = 07F;
    reg [9:0] I_filtered_10b[838] = 066;
    reg [9:0] I_filtered_10b[837] = 046;
    reg [9:0] I_filtered_10b[836] = 021;
    reg [9:0] I_filtered_10b[835] = 3F4;
    reg [9:0] I_filtered_10b[834] = 3C8;
    reg [9:0] I_filtered_10b[833] = 399;
    reg [9:0] I_filtered_10b[832] = 36D;
    reg [9:0] I_filtered_10b[831] = 349;
    reg [9:0] I_filtered_10b[830] = 32C;
    reg [9:0] I_filtered_10b[829] = 319;
    reg [9:0] I_filtered_10b[828] = 310;
    reg [9:0] I_filtered_10b[827] = 315;
    reg [9:0] I_filtered_10b[826] = 321;
    reg [9:0] I_filtered_10b[825] = 337;
    reg [9:0] I_filtered_10b[824] = 353;
    reg [9:0] I_filtered_10b[823] = 374;
    reg [9:0] I_filtered_10b[822] = 398;
    reg [9:0] I_filtered_10b[821] = 3B8;
    reg [9:0] I_filtered_10b[820] = 3D6;
    reg [9:0] I_filtered_10b[819] = 3EE;
    reg [9:0] I_filtered_10b[818] = 3FF;
    reg [9:0] I_filtered_10b[817] = 00E;
    reg [9:0] I_filtered_10b[816] = 01A;
    reg [9:0] I_filtered_10b[815] = 020;
    reg [9:0] I_filtered_10b[814] = 025;
    reg [9:0] I_filtered_10b[813] = 02F;
    reg [9:0] I_filtered_10b[812] = 039;
    reg [9:0] I_filtered_10b[811] = 042;
    reg [9:0] I_filtered_10b[810] = 053;
    reg [9:0] I_filtered_10b[809] = 066;
    reg [9:0] I_filtered_10b[808] = 07A;
    reg [9:0] I_filtered_10b[807] = 092;
    reg [9:0] I_filtered_10b[806] = 0A7;
    reg [9:0] I_filtered_10b[805] = 0BA;
    reg [9:0] I_filtered_10b[804] = 0C9;
    reg [9:0] I_filtered_10b[803] = 0D2;
    reg [9:0] I_filtered_10b[802] = 0D8;
    reg [9:0] I_filtered_10b[801] = 0D5;
    reg [9:0] I_filtered_10b[800] = 0CE;
    reg [9:0] I_filtered_10b[799] = 0BF;
    reg [9:0] I_filtered_10b[798] = 0AD;
    reg [9:0] I_filtered_10b[797] = 096;
    reg [9:0] I_filtered_10b[796] = 080;
    reg [9:0] I_filtered_10b[795] = 06B;
    reg [9:0] I_filtered_10b[794] = 054;
    reg [9:0] I_filtered_10b[793] = 043;
    reg [9:0] I_filtered_10b[792] = 034;
    reg [9:0] I_filtered_10b[791] = 028;
    reg [9:0] I_filtered_10b[790] = 01B;
    reg [9:0] I_filtered_10b[789] = 014;
    reg [9:0] I_filtered_10b[788] = 00B;
    reg [9:0] I_filtered_10b[787] = 003;
    reg [9:0] I_filtered_10b[786] = 3FD;
    reg [9:0] I_filtered_10b[785] = 3F7;
    reg [9:0] I_filtered_10b[784] = 3F0;
    reg [9:0] I_filtered_10b[783] = 3E7;
    reg [9:0] I_filtered_10b[782] = 3E2;
    reg [9:0] I_filtered_10b[781] = 3D8;
    reg [9:0] I_filtered_10b[780] = 3D1;
    reg [9:0] I_filtered_10b[779] = 3C9;
    reg [9:0] I_filtered_10b[778] = 3C3;
    reg [9:0] I_filtered_10b[777] = 3BB;
    reg [9:0] I_filtered_10b[776] = 3B3;
    reg [9:0] I_filtered_10b[775] = 3AD;
    reg [9:0] I_filtered_10b[774] = 3A3;
    reg [9:0] I_filtered_10b[773] = 39B;
    reg [9:0] I_filtered_10b[772] = 391;
    reg [9:0] I_filtered_10b[771] = 386;
    reg [9:0] I_filtered_10b[770] = 378;
    reg [9:0] I_filtered_10b[769] = 36C;
    reg [9:0] I_filtered_10b[768] = 35D;
    reg [9:0] I_filtered_10b[767] = 34E;
    reg [9:0] I_filtered_10b[766] = 340;
    reg [9:0] I_filtered_10b[765] = 336;
    reg [9:0] I_filtered_10b[764] = 330;
    reg [9:0] I_filtered_10b[763] = 32E;
    reg [9:0] I_filtered_10b[762] = 331;
    reg [9:0] I_filtered_10b[761] = 339;
    reg [9:0] I_filtered_10b[760] = 347;
    reg [9:0] I_filtered_10b[759] = 358;
    reg [9:0] I_filtered_10b[758] = 36D;
    reg [9:0] I_filtered_10b[757] = 386;
    reg [9:0] I_filtered_10b[756] = 39E;
    reg [9:0] I_filtered_10b[755] = 3B6;
    reg [9:0] I_filtered_10b[754] = 3CC;
    reg [9:0] I_filtered_10b[753] = 3DC;
    reg [9:0] I_filtered_10b[752] = 3E9;
    reg [9:0] I_filtered_10b[751] = 3F4;
    reg [9:0] I_filtered_10b[750] = 3F8;
    reg [9:0] I_filtered_10b[749] = 3F8;
    reg [9:0] I_filtered_10b[748] = 3F7;
    reg [9:0] I_filtered_10b[747] = 3F4;
    reg [9:0] I_filtered_10b[746] = 3F0;
    reg [9:0] I_filtered_10b[745] = 3EC;
    reg [9:0] I_filtered_10b[744] = 3E7;
    reg [9:0] I_filtered_10b[743] = 3E4;
    reg [9:0] I_filtered_10b[742] = 3E5;
    reg [9:0] I_filtered_10b[741] = 3E6;
    reg [9:0] I_filtered_10b[740] = 3EA;
    reg [9:0] I_filtered_10b[739] = 3EC;
    reg [9:0] I_filtered_10b[738] = 3EF;
    reg [9:0] I_filtered_10b[737] = 3F2;
    reg [9:0] I_filtered_10b[736] = 3F3;
    reg [9:0] I_filtered_10b[735] = 3EE;
    reg [9:0] I_filtered_10b[734] = 3E5;
    reg [9:0] I_filtered_10b[733] = 3DB;
    reg [9:0] I_filtered_10b[732] = 3CA;
    reg [9:0] I_filtered_10b[731] = 3B9;
    reg [9:0] I_filtered_10b[730] = 3A5;
    reg [9:0] I_filtered_10b[729] = 38F;
    reg [9:0] I_filtered_10b[728] = 37E;
    reg [9:0] I_filtered_10b[727] = 36E;
    reg [9:0] I_filtered_10b[726] = 362;
    reg [9:0] I_filtered_10b[725] = 35C;
    reg [9:0] I_filtered_10b[724] = 35B;
    reg [9:0] I_filtered_10b[723] = 360;
    reg [9:0] I_filtered_10b[722] = 36D;
    reg [9:0] I_filtered_10b[721] = 380;
    reg [9:0] I_filtered_10b[720] = 398;
    reg [9:0] I_filtered_10b[719] = 3B4;
    reg [9:0] I_filtered_10b[718] = 3D6;
    reg [9:0] I_filtered_10b[717] = 3F7;
    reg [9:0] I_filtered_10b[716] = 018;
    reg [9:0] I_filtered_10b[715] = 036;
    reg [9:0] I_filtered_10b[714] = 04D;
    reg [9:0] I_filtered_10b[713] = 061;
    reg [9:0] I_filtered_10b[712] = 06D;
    reg [9:0] I_filtered_10b[711] = 071;
    reg [9:0] I_filtered_10b[710] = 06E;
    reg [9:0] I_filtered_10b[709] = 067;
    reg [9:0] I_filtered_10b[708] = 05A;
    reg [9:0] I_filtered_10b[707] = 04A;
    reg [9:0] I_filtered_10b[706] = 039;
    reg [9:0] I_filtered_10b[705] = 026;
    reg [9:0] I_filtered_10b[704] = 016;
    reg [9:0] I_filtered_10b[703] = 008;
    reg [9:0] I_filtered_10b[702] = 3FD;
    reg [9:0] I_filtered_10b[701] = 3F5;
    reg [9:0] I_filtered_10b[700] = 3EE;
    reg [9:0] I_filtered_10b[699] = 3E8;
    reg [9:0] I_filtered_10b[698] = 3E6;
    reg [9:0] I_filtered_10b[697] = 3E3;
    reg [9:0] I_filtered_10b[696] = 3DD;
    reg [9:0] I_filtered_10b[695] = 3D6;
    reg [9:0] I_filtered_10b[694] = 3CF;
    reg [9:0] I_filtered_10b[693] = 3C2;
    reg [9:0] I_filtered_10b[692] = 3B6;
    reg [9:0] I_filtered_10b[691] = 3A8;
    reg [9:0] I_filtered_10b[690] = 397;
    reg [9:0] I_filtered_10b[689] = 38A;
    reg [9:0] I_filtered_10b[688] = 37D;
    reg [9:0] I_filtered_10b[687] = 373;
    reg [9:0] I_filtered_10b[686] = 36C;
    reg [9:0] I_filtered_10b[685] = 367;
    reg [9:0] I_filtered_10b[684] = 367;
    reg [9:0] I_filtered_10b[683] = 36B;
    reg [9:0] I_filtered_10b[682] = 375;
    reg [9:0] I_filtered_10b[681] = 381;
    reg [9:0] I_filtered_10b[680] = 391;
    reg [9:0] I_filtered_10b[679] = 3A2;
    reg [9:0] I_filtered_10b[678] = 3B4;
    reg [9:0] I_filtered_10b[677] = 3C7;
    reg [9:0] I_filtered_10b[676] = 3D6;
    reg [9:0] I_filtered_10b[675] = 3E3;
    reg [9:0] I_filtered_10b[674] = 3ED;
    reg [9:0] I_filtered_10b[673] = 3F5;
    reg [9:0] I_filtered_10b[672] = 3F8;
    reg [9:0] I_filtered_10b[671] = 3F9;
    reg [9:0] I_filtered_10b[670] = 3F5;
    reg [9:0] I_filtered_10b[669] = 3EF;
    reg [9:0] I_filtered_10b[668] = 3E6;
    reg [9:0] I_filtered_10b[667] = 3DB;
    reg [9:0] I_filtered_10b[666] = 3CF;
    reg [9:0] I_filtered_10b[665] = 3C2;
    reg [9:0] I_filtered_10b[664] = 3B7;
    reg [9:0] I_filtered_10b[663] = 3AD;
    reg [9:0] I_filtered_10b[662] = 3A6;
    reg [9:0] I_filtered_10b[661] = 3A0;
    reg [9:0] I_filtered_10b[660] = 39F;
    reg [9:0] I_filtered_10b[659] = 3A1;
    reg [9:0] I_filtered_10b[658] = 3A5;
    reg [9:0] I_filtered_10b[657] = 3AD;
    reg [9:0] I_filtered_10b[656] = 3B6;
    reg [9:0] I_filtered_10b[655] = 3C3;
    reg [9:0] I_filtered_10b[654] = 3D0;
    reg [9:0] I_filtered_10b[653] = 3E1;
    reg [9:0] I_filtered_10b[652] = 3EF;
    reg [9:0] I_filtered_10b[651] = 3FD;
    reg [9:0] I_filtered_10b[650] = 00B;
    reg [9:0] I_filtered_10b[649] = 015;
    reg [9:0] I_filtered_10b[648] = 01E;
    reg [9:0] I_filtered_10b[647] = 023;
    reg [9:0] I_filtered_10b[646] = 026;
    reg [9:0] I_filtered_10b[645] = 024;
    reg [9:0] I_filtered_10b[644] = 024;
    reg [9:0] I_filtered_10b[643] = 022;
    reg [9:0] I_filtered_10b[642] = 01F;
    reg [9:0] I_filtered_10b[641] = 01E;
    reg [9:0] I_filtered_10b[640] = 01C;
    reg [9:0] I_filtered_10b[639] = 01D;
    reg [9:0] I_filtered_10b[638] = 020;
    reg [9:0] I_filtered_10b[637] = 023;
    reg [9:0] I_filtered_10b[636] = 028;
    reg [9:0] I_filtered_10b[635] = 02B;
    reg [9:0] I_filtered_10b[634] = 02B;
    reg [9:0] I_filtered_10b[633] = 02C;
    reg [9:0] I_filtered_10b[632] = 028;
    reg [9:0] I_filtered_10b[631] = 01F;
    reg [9:0] I_filtered_10b[630] = 012;
    reg [9:0] I_filtered_10b[629] = 002;
    reg [9:0] I_filtered_10b[628] = 3ED;
    reg [9:0] I_filtered_10b[627] = 3D4;
    reg [9:0] I_filtered_10b[626] = 3B9;
    reg [9:0] I_filtered_10b[625] = 39F;
    reg [9:0] I_filtered_10b[624] = 386;
    reg [9:0] I_filtered_10b[623] = 374;
    reg [9:0] I_filtered_10b[622] = 365;
    reg [9:0] I_filtered_10b[621] = 35D;
    reg [9:0] I_filtered_10b[620] = 35B;
    reg [9:0] I_filtered_10b[619] = 362;
    reg [9:0] I_filtered_10b[618] = 36C;
    reg [9:0] I_filtered_10b[617] = 37C;
    reg [9:0] I_filtered_10b[616] = 38F;
    reg [9:0] I_filtered_10b[615] = 3A5;
    reg [9:0] I_filtered_10b[614] = 3BD;
    reg [9:0] I_filtered_10b[613] = 3D1;
    reg [9:0] I_filtered_10b[612] = 3E5;
    reg [9:0] I_filtered_10b[611] = 3F5;
    reg [9:0] I_filtered_10b[610] = 000;
    reg [9:0] I_filtered_10b[609] = 00B;
    reg [9:0] I_filtered_10b[608] = 014;
    reg [9:0] I_filtered_10b[607] = 01A;
    reg [9:0] I_filtered_10b[606] = 01F;
    reg [9:0] I_filtered_10b[605] = 029;
    reg [9:0] I_filtered_10b[604] = 034;
    reg [9:0] I_filtered_10b[603] = 040;
    reg [9:0] I_filtered_10b[602] = 051;
    reg [9:0] I_filtered_10b[601] = 064;
    reg [9:0] I_filtered_10b[600] = 077;
    reg [9:0] I_filtered_10b[599] = 091;
    reg [9:0] I_filtered_10b[598] = 0A5;
    reg [9:0] I_filtered_10b[597] = 0BC;
    reg [9:0] I_filtered_10b[596] = 0CC;
    reg [9:0] I_filtered_10b[595] = 0D7;
    reg [9:0] I_filtered_10b[594] = 0DE;
    reg [9:0] I_filtered_10b[593] = 0DE;
    reg [9:0] I_filtered_10b[592] = 0D5;
    reg [9:0] I_filtered_10b[591] = 0C2;
    reg [9:0] I_filtered_10b[590] = 0AA;
    reg [9:0] I_filtered_10b[589] = 08A;
    reg [9:0] I_filtered_10b[588] = 069;
    reg [9:0] I_filtered_10b[587] = 045;
    reg [9:0] I_filtered_10b[586] = 01F;
    reg [9:0] I_filtered_10b[585] = 000;
    reg [9:0] I_filtered_10b[584] = 3E2;
    reg [9:0] I_filtered_10b[583] = 3CC;
    reg [9:0] I_filtered_10b[582] = 3BD;
    reg [9:0] I_filtered_10b[581] = 3B6;
    reg [9:0] I_filtered_10b[580] = 3B7;
    reg [9:0] I_filtered_10b[579] = 3C2;
    reg [9:0] I_filtered_10b[578] = 3D8;
    reg [9:0] I_filtered_10b[577] = 3F4;
    reg [9:0] I_filtered_10b[576] = 017;
    reg [9:0] I_filtered_10b[575] = 03D;
    reg [9:0] I_filtered_10b[574] = 067;
    reg [9:0] I_filtered_10b[573] = 090;
    reg [9:0] I_filtered_10b[572] = 0B4;
    reg [9:0] I_filtered_10b[571] = 0D4;
    reg [9:0] I_filtered_10b[570] = 0EB;
    reg [9:0] I_filtered_10b[569] = 0F6;
    reg [9:0] I_filtered_10b[568] = 0F6;
    reg [9:0] I_filtered_10b[567] = 0ED;
    reg [9:0] I_filtered_10b[566] = 0D6;
    reg [9:0] I_filtered_10b[565] = 0B4;
    reg [9:0] I_filtered_10b[564] = 087;
    reg [9:0] I_filtered_10b[563] = 055;
    reg [9:0] I_filtered_10b[562] = 019;
    reg [9:0] I_filtered_10b[561] = 3E0;
    reg [9:0] I_filtered_10b[560] = 3A6;
    reg [9:0] I_filtered_10b[559] = 370;
    reg [9:0] I_filtered_10b[558] = 344;
    reg [9:0] I_filtered_10b[557] = 321;
    reg [9:0] I_filtered_10b[556] = 30B;
    reg [9:0] I_filtered_10b[555] = 304;
    reg [9:0] I_filtered_10b[554] = 309;
    reg [9:0] I_filtered_10b[553] = 319;
    reg [9:0] I_filtered_10b[552] = 335;
    reg [9:0] I_filtered_10b[551] = 359;
    reg [9:0] I_filtered_10b[550] = 383;
    reg [9:0] I_filtered_10b[549] = 3B2;
    reg [9:0] I_filtered_10b[548] = 3DE;
    reg [9:0] I_filtered_10b[547] = 007;
    reg [9:0] I_filtered_10b[546] = 02C;
    reg [9:0] I_filtered_10b[545] = 048;
    reg [9:0] I_filtered_10b[544] = 05F;
    reg [9:0] I_filtered_10b[543] = 06E;
    reg [9:0] I_filtered_10b[542] = 071;
    reg [9:0] I_filtered_10b[541] = 070;
    reg [9:0] I_filtered_10b[540] = 06B;
    reg [9:0] I_filtered_10b[539] = 062;
    reg [9:0] I_filtered_10b[538] = 054;
    reg [9:0] I_filtered_10b[537] = 049;
    reg [9:0] I_filtered_10b[536] = 03D;
    reg [9:0] I_filtered_10b[535] = 033;
    reg [9:0] I_filtered_10b[534] = 02C;
    reg [9:0] I_filtered_10b[533] = 026;
    reg [9:0] I_filtered_10b[532] = 020;
    reg [9:0] I_filtered_10b[531] = 01D;
    reg [9:0] I_filtered_10b[530] = 019;
    reg [9:0] I_filtered_10b[529] = 01A;
    reg [9:0] I_filtered_10b[528] = 017;
    reg [9:0] I_filtered_10b[527] = 014;
    reg [9:0] I_filtered_10b[526] = 011;
    reg [9:0] I_filtered_10b[525] = 00F;
    reg [9:0] I_filtered_10b[524] = 009;
    reg [9:0] I_filtered_10b[523] = 004;
    reg [9:0] I_filtered_10b[522] = 000;
    reg [9:0] I_filtered_10b[521] = 3FB;
    reg [9:0] I_filtered_10b[520] = 3F8;
    reg [9:0] I_filtered_10b[519] = 3F6;
    reg [9:0] I_filtered_10b[518] = 3F4;
    reg [9:0] I_filtered_10b[517] = 3F0;
    reg [9:0] I_filtered_10b[516] = 3EC;
    reg [9:0] I_filtered_10b[515] = 3E9;
    reg [9:0] I_filtered_10b[514] = 3E1;
    reg [9:0] I_filtered_10b[513] = 3D9;
    reg [9:0] I_filtered_10b[512] = 3CE;
    reg [9:0] I_filtered_10b[511] = 3C2;
    reg [9:0] I_filtered_10b[510] = 3B4;
    reg [9:0] I_filtered_10b[509] = 3A6;
    reg [9:0] I_filtered_10b[508] = 395;
    reg [9:0] I_filtered_10b[507] = 386;
    reg [9:0] I_filtered_10b[506] = 377;
    reg [9:0] I_filtered_10b[505] = 36C;
    reg [9:0] I_filtered_10b[504] = 365;
    reg [9:0] I_filtered_10b[503] = 361;
    reg [9:0] I_filtered_10b[502] = 362;
    reg [9:0] I_filtered_10b[501] = 36A;
    reg [9:0] I_filtered_10b[500] = 378;
    reg [9:0] I_filtered_10b[499] = 38A;
    reg [9:0] I_filtered_10b[498] = 3A1;
    reg [9:0] I_filtered_10b[497] = 3BA;
    reg [9:0] I_filtered_10b[496] = 3D4;
    reg [9:0] I_filtered_10b[495] = 3F0;
    reg [9:0] I_filtered_10b[494] = 007;
    reg [9:0] I_filtered_10b[493] = 01D;
    reg [9:0] I_filtered_10b[492] = 02D;
    reg [9:0] I_filtered_10b[491] = 039;
    reg [9:0] I_filtered_10b[490] = 03E;
    reg [9:0] I_filtered_10b[489] = 03D;
    reg [9:0] I_filtered_10b[488] = 035;
    reg [9:0] I_filtered_10b[487] = 024;
    reg [9:0] I_filtered_10b[486] = 010;
    reg [9:0] I_filtered_10b[485] = 3F6;
    reg [9:0] I_filtered_10b[484] = 3D7;
    reg [9:0] I_filtered_10b[483] = 3B5;
    reg [9:0] I_filtered_10b[482] = 397;
    reg [9:0] I_filtered_10b[481] = 37A;
    reg [9:0] I_filtered_10b[480] = 365;
    reg [9:0] I_filtered_10b[479] = 353;
    reg [9:0] I_filtered_10b[478] = 34D;
    reg [9:0] I_filtered_10b[477] = 34F;
    reg [9:0] I_filtered_10b[476] = 35A;
    reg [9:0] I_filtered_10b[475] = 36D;
    reg [9:0] I_filtered_10b[474] = 386;
    reg [9:0] I_filtered_10b[473] = 3A6;
    reg [9:0] I_filtered_10b[472] = 3C8;
    reg [9:0] I_filtered_10b[471] = 3EF;
    reg [9:0] I_filtered_10b[470] = 00F;
    reg [9:0] I_filtered_10b[469] = 032;
    reg [9:0] I_filtered_10b[468] = 050;
    reg [9:0] I_filtered_10b[467] = 06A;
    reg [9:0] I_filtered_10b[466] = 07F;
    reg [9:0] I_filtered_10b[465] = 090;
    reg [9:0] I_filtered_10b[464] = 099;
    reg [9:0] I_filtered_10b[463] = 09F;
    reg [9:0] I_filtered_10b[462] = 0A5;
    reg [9:0] I_filtered_10b[461] = 0A5;
    reg [9:0] I_filtered_10b[460] = 0A4;
    reg [9:0] I_filtered_10b[459] = 0A5;
    reg [9:0] I_filtered_10b[458] = 0A6;
    reg [9:0] I_filtered_10b[457] = 0A6;
    reg [9:0] I_filtered_10b[456] = 0AB;
    reg [9:0] I_filtered_10b[455] = 0AE;
    reg [9:0] I_filtered_10b[454] = 0B4;
    reg [9:0] I_filtered_10b[453] = 0B8;
    reg [9:0] I_filtered_10b[452] = 0BC;
    reg [9:0] I_filtered_10b[451] = 0C0;
    reg [9:0] I_filtered_10b[450] = 0C2;
    reg [9:0] I_filtered_10b[449] = 0C2;
    reg [9:0] I_filtered_10b[448] = 0BE;
    reg [9:0] I_filtered_10b[447] = 0BA;
    reg [9:0] I_filtered_10b[446] = 0B3;
    reg [9:0] I_filtered_10b[445] = 0AE;
    reg [9:0] I_filtered_10b[444] = 0A7;
    reg [9:0] I_filtered_10b[443] = 09E;
    reg [9:0] I_filtered_10b[442] = 099;
    reg [9:0] I_filtered_10b[441] = 092;
    reg [9:0] I_filtered_10b[440] = 08E;
    reg [9:0] I_filtered_10b[439] = 086;
    reg [9:0] I_filtered_10b[438] = 081;
    reg [9:0] I_filtered_10b[437] = 07B;
    reg [9:0] I_filtered_10b[436] = 076;
    reg [9:0] I_filtered_10b[435] = 074;
    reg [9:0] I_filtered_10b[434] = 070;
    reg [9:0] I_filtered_10b[433] = 06F;
    reg [9:0] I_filtered_10b[432] = 06B;
    reg [9:0] I_filtered_10b[431] = 06C;
    reg [9:0] I_filtered_10b[430] = 06C;
    reg [9:0] I_filtered_10b[429] = 06A;
    reg [9:0] I_filtered_10b[428] = 06B;
    reg [9:0] I_filtered_10b[427] = 06A;
    reg [9:0] I_filtered_10b[426] = 065;
    reg [9:0] I_filtered_10b[425] = 05F;
    reg [9:0] I_filtered_10b[424] = 059;
    reg [9:0] I_filtered_10b[423] = 04C;
    reg [9:0] I_filtered_10b[422] = 03B;
    reg [9:0] I_filtered_10b[421] = 026;
    reg [9:0] I_filtered_10b[420] = 00D;
    reg [9:0] I_filtered_10b[419] = 3EF;
    reg [9:0] I_filtered_10b[418] = 3D0;
    reg [9:0] I_filtered_10b[417] = 3AE;
    reg [9:0] I_filtered_10b[416] = 38D;
    reg [9:0] I_filtered_10b[415] = 372;
    reg [9:0] I_filtered_10b[414] = 35C;
    reg [9:0] I_filtered_10b[413] = 34F;
    reg [9:0] I_filtered_10b[412] = 349;
    reg [9:0] I_filtered_10b[411] = 34F;
    reg [9:0] I_filtered_10b[410] = 35F;
    reg [9:0] I_filtered_10b[409] = 378;
    reg [9:0] I_filtered_10b[408] = 397;
    reg [9:0] I_filtered_10b[407] = 3BE;
    reg [9:0] I_filtered_10b[406] = 3EA;
    reg [9:0] I_filtered_10b[405] = 014;
    reg [9:0] I_filtered_10b[404] = 03D;
    reg [9:0] I_filtered_10b[403] = 061;
    reg [9:0] I_filtered_10b[402] = 07C;
    reg [9:0] I_filtered_10b[401] = 092;
    reg [9:0] I_filtered_10b[400] = 0A0;
    reg [9:0] I_filtered_10b[399] = 0A5;
    reg [9:0] I_filtered_10b[398] = 0A2;
    reg [9:0] I_filtered_10b[397] = 09E;
    reg [9:0] I_filtered_10b[396] = 096;
    reg [9:0] I_filtered_10b[395] = 089;
    reg [9:0] I_filtered_10b[394] = 07F;
    reg [9:0] I_filtered_10b[393] = 073;
    reg [9:0] I_filtered_10b[392] = 06C;
    reg [9:0] I_filtered_10b[391] = 068;
    reg [9:0] I_filtered_10b[390] = 064;
    reg [9:0] I_filtered_10b[389] = 064;
    reg [9:0] I_filtered_10b[388] = 063;
    reg [9:0] I_filtered_10b[387] = 060;
    reg [9:0] I_filtered_10b[386] = 05F;
    reg [9:0] I_filtered_10b[385] = 05A;
    reg [9:0] I_filtered_10b[384] = 04F;
    reg [9:0] I_filtered_10b[383] = 03E;
    reg [9:0] I_filtered_10b[382] = 02C;
    reg [9:0] I_filtered_10b[381] = 011;
    reg [9:0] I_filtered_10b[380] = 3F6;
    reg [9:0] I_filtered_10b[379] = 3DA;
    reg [9:0] I_filtered_10b[378] = 3B8;
    reg [9:0] I_filtered_10b[377] = 39D;
    reg [9:0] I_filtered_10b[376] = 382;
    reg [9:0] I_filtered_10b[375] = 36E;
    reg [9:0] I_filtered_10b[374] = 35E;
    reg [9:0] I_filtered_10b[373] = 355;
    reg [9:0] I_filtered_10b[372] = 353;
    reg [9:0] I_filtered_10b[371] = 359;
    reg [9:0] I_filtered_10b[370] = 36A;
    reg [9:0] I_filtered_10b[369] = 37E;
    reg [9:0] I_filtered_10b[368] = 399;
    reg [9:0] I_filtered_10b[367] = 3B5;
    reg [9:0] I_filtered_10b[366] = 3D5;
    reg [9:0] I_filtered_10b[365] = 3F4;
    reg [9:0] I_filtered_10b[364] = 00E;
    reg [9:0] I_filtered_10b[363] = 025;
    reg [9:0] I_filtered_10b[362] = 037;
    reg [9:0] I_filtered_10b[361] = 041;
    reg [9:0] I_filtered_10b[360] = 044;
    reg [9:0] I_filtered_10b[359] = 041;
    reg [9:0] I_filtered_10b[358] = 034;
    reg [9:0] I_filtered_10b[357] = 01F;
    reg [9:0] I_filtered_10b[356] = 004;
    reg [9:0] I_filtered_10b[355] = 3E4;
    reg [9:0] I_filtered_10b[354] = 3C0;
    reg [9:0] I_filtered_10b[353] = 39A;
    reg [9:0] I_filtered_10b[352] = 374;
    reg [9:0] I_filtered_10b[351] = 353;
    reg [9:0] I_filtered_10b[350] = 334;
    reg [9:0] I_filtered_10b[349] = 31E;
    reg [9:0] I_filtered_10b[348] = 312;
    reg [9:0] I_filtered_10b[347] = 310;
    reg [9:0] I_filtered_10b[346] = 316;
    reg [9:0] I_filtered_10b[345] = 329;
    reg [9:0] I_filtered_10b[344] = 346;
    reg [9:0] I_filtered_10b[343] = 36D;
    reg [9:0] I_filtered_10b[342] = 399;
    reg [9:0] I_filtered_10b[341] = 3CE;
    reg [9:0] I_filtered_10b[340] = 002;
    reg [9:0] I_filtered_10b[339] = 036;
    reg [9:0] I_filtered_10b[338] = 067;
    reg [9:0] I_filtered_10b[337] = 08D;
    reg [9:0] I_filtered_10b[336] = 0AC;
    reg [9:0] I_filtered_10b[335] = 0BE;
    reg [9:0] I_filtered_10b[334] = 0C3;
    reg [9:0] I_filtered_10b[333] = 0BB;
    reg [9:0] I_filtered_10b[332] = 0AA;
    reg [9:0] I_filtered_10b[331] = 08E;
    reg [9:0] I_filtered_10b[330] = 06B;
    reg [9:0] I_filtered_10b[329] = 043;
    reg [9:0] I_filtered_10b[328] = 017;
    reg [9:0] I_filtered_10b[327] = 3EF;
    reg [9:0] I_filtered_10b[326] = 3C8;
    reg [9:0] I_filtered_10b[325] = 3A7;
    reg [9:0] I_filtered_10b[324] = 38C;
    reg [9:0] I_filtered_10b[323] = 376;
    reg [9:0] I_filtered_10b[322] = 367;
    reg [9:0] I_filtered_10b[321] = 361;
    reg [9:0] I_filtered_10b[320] = 35E;
    reg [9:0] I_filtered_10b[319] = 35D;
    reg [9:0] I_filtered_10b[318] = 361;
    reg [9:0] I_filtered_10b[317] = 369;
    reg [9:0] I_filtered_10b[316] = 36E;
    reg [9:0] I_filtered_10b[315] = 373;
    reg [9:0] I_filtered_10b[314] = 378;
    reg [9:0] I_filtered_10b[313] = 37A;
    reg [9:0] I_filtered_10b[312] = 37D;
    reg [9:0] I_filtered_10b[311] = 37F;
    reg [9:0] I_filtered_10b[310] = 380;
    reg [9:0] I_filtered_10b[309] = 381;
    reg [9:0] I_filtered_10b[308] = 37F;
    reg [9:0] I_filtered_10b[307] = 380;
    reg [9:0] I_filtered_10b[306] = 37E;
    reg [9:0] I_filtered_10b[305] = 37D;
    reg [9:0] I_filtered_10b[304] = 37A;
    reg [9:0] I_filtered_10b[303] = 378;
    reg [9:0] I_filtered_10b[302] = 376;
    reg [9:0] I_filtered_10b[301] = 372;
    reg [9:0] I_filtered_10b[300] = 36E;
    reg [9:0] I_filtered_10b[299] = 36A;
    reg [9:0] I_filtered_10b[298] = 365;
    reg [9:0] I_filtered_10b[297] = 362;
    reg [9:0] I_filtered_10b[296] = 364;
    reg [9:0] I_filtered_10b[295] = 367;
    reg [9:0] I_filtered_10b[294] = 36D;
    reg [9:0] I_filtered_10b[293] = 37A;
    reg [9:0] I_filtered_10b[292] = 38B;
    reg [9:0] I_filtered_10b[291] = 3A1;
    reg [9:0] I_filtered_10b[290] = 3BA;
    reg [9:0] I_filtered_10b[289] = 3D7;
    reg [9:0] I_filtered_10b[288] = 3F2;
    reg [9:0] I_filtered_10b[287] = 012;
    reg [9:0] I_filtered_10b[286] = 02E;
    reg [9:0] I_filtered_10b[285] = 04A;
    reg [9:0] I_filtered_10b[284] = 05E;
    reg [9:0] I_filtered_10b[283] = 06E;
    reg [9:0] I_filtered_10b[282] = 077;
    reg [9:0] I_filtered_10b[281] = 079;
    reg [9:0] I_filtered_10b[280] = 073;
    reg [9:0] I_filtered_10b[279] = 062;
    reg [9:0] I_filtered_10b[278] = 04D;
    reg [9:0] I_filtered_10b[277] = 031;
    reg [9:0] I_filtered_10b[276] = 013;
    reg [9:0] I_filtered_10b[275] = 3F1;
    reg [9:0] I_filtered_10b[274] = 3D1;
    reg [9:0] I_filtered_10b[273] = 3B5;
    reg [9:0] I_filtered_10b[272] = 39D;
    reg [9:0] I_filtered_10b[271] = 38B;
    reg [9:0] I_filtered_10b[270] = 383;
    reg [9:0] I_filtered_10b[269] = 383;
    reg [9:0] I_filtered_10b[268] = 38A;
    reg [9:0] I_filtered_10b[267] = 39B;
    reg [9:0] I_filtered_10b[266] = 3B4;
    reg [9:0] I_filtered_10b[265] = 3D5;
    reg [9:0] I_filtered_10b[264] = 3FA;
    reg [9:0] I_filtered_10b[263] = 023;
    reg [9:0] I_filtered_10b[262] = 04B;
    reg [9:0] I_filtered_10b[261] = 075;
    reg [9:0] I_filtered_10b[260] = 099;
    reg [9:0] I_filtered_10b[259] = 0BB;
    reg [9:0] I_filtered_10b[258] = 0D4;
    reg [9:0] I_filtered_10b[257] = 0E4;
    reg [9:0] I_filtered_10b[256] = 0EA;
    reg [9:0] I_filtered_10b[255] = 0E9;
    reg [9:0] I_filtered_10b[254] = 0DE;
    reg [9:0] I_filtered_10b[253] = 0C9;
    reg [9:0] I_filtered_10b[252] = 0AC;
    reg [9:0] I_filtered_10b[251] = 08B;
    reg [9:0] I_filtered_10b[250] = 066;
    reg [9:0] I_filtered_10b[249] = 040;
    reg [9:0] I_filtered_10b[248] = 01B;
    reg [9:0] I_filtered_10b[247] = 3FA;
    reg [9:0] I_filtered_10b[246] = 3DD;
    reg [9:0] I_filtered_10b[245] = 3C7;
    reg [9:0] I_filtered_10b[244] = 3BA;
    reg [9:0] I_filtered_10b[243] = 3B6;
    reg [9:0] I_filtered_10b[242] = 3BA;
    reg [9:0] I_filtered_10b[241] = 3C7;
    reg [9:0] I_filtered_10b[240] = 3DD;
    reg [9:0] I_filtered_10b[239] = 3FA;
    reg [9:0] I_filtered_10b[238] = 01B;
    reg [9:0] I_filtered_10b[237] = 041;
    reg [9:0] I_filtered_10b[236] = 068;
    reg [9:0] I_filtered_10b[235] = 08D;
    reg [9:0] I_filtered_10b[234] = 0AF;
    reg [9:0] I_filtered_10b[233] = 0CB;
    reg [9:0] I_filtered_10b[232] = 0E0;
    reg [9:0] I_filtered_10b[231] = 0EA;
    reg [9:0] I_filtered_10b[230] = 0EA;
    reg [9:0] I_filtered_10b[229] = 0E2;
    reg [9:0] I_filtered_10b[228] = 0D1;
    reg [9:0] I_filtered_10b[227] = 0B8;
    reg [9:0] I_filtered_10b[226] = 096;
    reg [9:0] I_filtered_10b[225] = 073;
    reg [9:0] I_filtered_10b[224] = 04A;
    reg [9:0] I_filtered_10b[223] = 025;
    reg [9:0] I_filtered_10b[222] = 3FF;
    reg [9:0] I_filtered_10b[221] = 3DD;
    reg [9:0] I_filtered_10b[220] = 3BF;
    reg [9:0] I_filtered_10b[219] = 3A8;
    reg [9:0] I_filtered_10b[218] = 397;
    reg [9:0] I_filtered_10b[217] = 38F;
    reg [9:0] I_filtered_10b[216] = 38C;
    reg [9:0] I_filtered_10b[215] = 38D;
    reg [9:0] I_filtered_10b[214] = 396;
    reg [9:0] I_filtered_10b[213] = 3A3;
    reg [9:0] I_filtered_10b[212] = 3B1;
    reg [9:0] I_filtered_10b[211] = 3BF;
    reg [9:0] I_filtered_10b[210] = 3CF;
    reg [9:0] I_filtered_10b[209] = 3DC;
    reg [9:0] I_filtered_10b[208] = 3E8;
    reg [9:0] I_filtered_10b[207] = 3F1;
    reg [9:0] I_filtered_10b[206] = 3F8;
    reg [9:0] I_filtered_10b[205] = 3FB;
    reg [9:0] I_filtered_10b[204] = 3F8;
    reg [9:0] I_filtered_10b[203] = 3F6;
    reg [9:0] I_filtered_10b[202] = 3ED;
    reg [9:0] I_filtered_10b[201] = 3E3;
    reg [9:0] I_filtered_10b[200] = 3D5;
    reg [9:0] I_filtered_10b[199] = 3C6;
    reg [9:0] I_filtered_10b[198] = 3B5;
    reg [9:0] I_filtered_10b[197] = 3A4;
    reg [9:0] I_filtered_10b[196] = 391;
    reg [9:0] I_filtered_10b[195] = 381;
    reg [9:0] I_filtered_10b[194] = 36F;
    reg [9:0] I_filtered_10b[193] = 363;
    reg [9:0] I_filtered_10b[192] = 35D;
    reg [9:0] I_filtered_10b[191] = 35B;
    reg [9:0] I_filtered_10b[190] = 35E;
    reg [9:0] I_filtered_10b[189] = 369;
    reg [9:0] I_filtered_10b[188] = 37C;
    reg [9:0] I_filtered_10b[187] = 395;
    reg [9:0] I_filtered_10b[186] = 3B2;
    reg [9:0] I_filtered_10b[185] = 3D6;
    reg [9:0] I_filtered_10b[184] = 3FC;
    reg [9:0] I_filtered_10b[183] = 020;
    reg [9:0] I_filtered_10b[182] = 044;
    reg [9:0] I_filtered_10b[181] = 05F;
    reg [9:0] I_filtered_10b[180] = 075;
    reg [9:0] I_filtered_10b[179] = 081;
    reg [9:0] I_filtered_10b[178] = 083;
    reg [9:0] I_filtered_10b[177] = 07A;
    reg [9:0] I_filtered_10b[176] = 068;
    reg [9:0] I_filtered_10b[175] = 04E;
    reg [9:0] I_filtered_10b[174] = 02E;
    reg [9:0] I_filtered_10b[173] = 008;
    reg [9:0] I_filtered_10b[172] = 3DF;
    reg [9:0] I_filtered_10b[171] = 3BA;
    reg [9:0] I_filtered_10b[170] = 394;
    reg [9:0] I_filtered_10b[169] = 375;
    reg [9:0] I_filtered_10b[168] = 35A;
    reg [9:0] I_filtered_10b[167] = 345;
    reg [9:0] I_filtered_10b[166] = 335;
    reg [9:0] I_filtered_10b[165] = 32E;
    reg [9:0] I_filtered_10b[164] = 329;
    reg [9:0] I_filtered_10b[163] = 327;
    reg [9:0] I_filtered_10b[162] = 32A;
    reg [9:0] I_filtered_10b[161] = 331;
    reg [9:0] I_filtered_10b[160] = 336;
    reg [9:0] I_filtered_10b[159] = 33A;
    reg [9:0] I_filtered_10b[158] = 33E;
    reg [9:0] I_filtered_10b[157] = 341;
    reg [9:0] I_filtered_10b[156] = 344;
    reg [9:0] I_filtered_10b[155] = 347;
    reg [9:0] I_filtered_10b[154] = 349;
    reg [9:0] I_filtered_10b[153] = 34C;
    reg [9:0] I_filtered_10b[152] = 34C;
    reg [9:0] I_filtered_10b[151] = 34F;
    reg [9:0] I_filtered_10b[150] = 34E;
    reg [9:0] I_filtered_10b[149] = 34C;
    reg [9:0] I_filtered_10b[148] = 34A;
    reg [9:0] I_filtered_10b[147] = 345;
    reg [9:0] I_filtered_10b[146] = 33F;
    reg [9:0] I_filtered_10b[145] = 334;
    reg [9:0] I_filtered_10b[144] = 32C;
    reg [9:0] I_filtered_10b[143] = 322;
    reg [9:0] I_filtered_10b[142] = 31A;
    reg [9:0] I_filtered_10b[141] = 315;
    reg [9:0] I_filtered_10b[140] = 31A;
    reg [9:0] I_filtered_10b[139] = 322;
    reg [9:0] I_filtered_10b[138] = 331;
    reg [9:0] I_filtered_10b[137] = 34A;
    reg [9:0] I_filtered_10b[136] = 368;
    reg [9:0] I_filtered_10b[135] = 38F;
    reg [9:0] I_filtered_10b[134] = 3B9;
    reg [9:0] I_filtered_10b[133] = 3EB;
    reg [9:0] I_filtered_10b[132] = 016;
    reg [9:0] I_filtered_10b[131] = 048;
    reg [9:0] I_filtered_10b[130] = 074;
    reg [9:0] I_filtered_10b[129] = 09C;
    reg [9:0] I_filtered_10b[128] = 0BB;
    reg [9:0] I_filtered_10b[127] = 0D5;
    reg [9:0] I_filtered_10b[126] = 0E4;
    reg [9:0] I_filtered_10b[125] = 0EB;
    reg [9:0] I_filtered_10b[124] = 0ED;
    reg [9:0] I_filtered_10b[123] = 0E3;
    reg [9:0] I_filtered_10b[122] = 0D7;
    reg [9:0] I_filtered_10b[121] = 0C5;
    reg [9:0] I_filtered_10b[120] = 0B6;
    reg [9:0] I_filtered_10b[119] = 0A3;
    reg [9:0] I_filtered_10b[118] = 093;
    reg [9:0] I_filtered_10b[117] = 088;
    reg [9:0] I_filtered_10b[116] = 07E;
    reg [9:0] I_filtered_10b[115] = 078;
    reg [9:0] I_filtered_10b[114] = 073;
    reg [9:0] I_filtered_10b[113] = 075;
    reg [9:0] I_filtered_10b[112] = 075;
    reg [9:0] I_filtered_10b[111] = 07A;
    reg [9:0] I_filtered_10b[110] = 081;
    reg [9:0] I_filtered_10b[109] = 08B;
    reg [9:0] I_filtered_10b[108] = 095;
    reg [9:0] I_filtered_10b[107] = 0A2;
    reg [9:0] I_filtered_10b[106] = 0B0;
    reg [9:0] I_filtered_10b[105] = 0BE;
    reg [9:0] I_filtered_10b[104] = 0CB;
    reg [9:0] I_filtered_10b[103] = 0D9;
    reg [9:0] I_filtered_10b[102] = 0E2;
    reg [9:0] I_filtered_10b[101] = 0E2;
    reg [9:0] I_filtered_10b[100] = 0DE;
    reg [9:0] I_filtered_10b[99] = 0D5;
    reg [9:0] I_filtered_10b[98] = 0C1;
    reg [9:0] I_filtered_10b[97] = 0A7;
    reg [9:0] I_filtered_10b[96] = 084;
    reg [9:0] I_filtered_10b[95] = 05D;
    reg [9:0] I_filtered_10b[94] = 02E;
    reg [9:0] I_filtered_10b[93] = 001;
    reg [9:0] I_filtered_10b[92] = 3D1;
    reg [9:0] I_filtered_10b[91] = 3A5;
    reg [9:0] I_filtered_10b[90] = 37F;
    reg [9:0] I_filtered_10b[89] = 361;
    reg [9:0] I_filtered_10b[88] = 34D;
    reg [9:0] I_filtered_10b[87] = 343;
    reg [9:0] I_filtered_10b[86] = 346;
    reg [9:0] I_filtered_10b[85] = 351;
    reg [9:0] I_filtered_10b[84] = 368;
    reg [9:0] I_filtered_10b[83] = 385;
    reg [9:0] I_filtered_10b[82] = 3A8;
    reg [9:0] I_filtered_10b[81] = 3CE;
    reg [9:0] I_filtered_10b[80] = 3F4;
    reg [9:0] I_filtered_10b[79] = 016;
    reg [9:0] I_filtered_10b[78] = 034;
    reg [9:0] I_filtered_10b[77] = 04B;
    reg [9:0] I_filtered_10b[76] = 05D;
    reg [9:0] I_filtered_10b[75] = 069;
    reg [9:0] I_filtered_10b[74] = 06B;
    reg [9:0] I_filtered_10b[73] = 06A;
    reg [9:0] I_filtered_10b[72] = 066;
    reg [9:0] I_filtered_10b[71] = 05E;
    reg [9:0] I_filtered_10b[70] = 052;
    reg [9:0] I_filtered_10b[69] = 048;
    reg [9:0] I_filtered_10b[68] = 03C;
    reg [9:0] I_filtered_10b[67] = 033;
    reg [9:0] I_filtered_10b[66] = 02B;
    reg [9:0] I_filtered_10b[65] = 023;
    reg [9:0] I_filtered_10b[64] = 01C;
    reg [9:0] I_filtered_10b[63] = 018;
    reg [9:0] I_filtered_10b[62] = 014;
    reg [9:0] I_filtered_10b[61] = 014;
    reg [9:0] I_filtered_10b[60] = 012;
    reg [9:0] I_filtered_10b[59] = 012;
    reg [9:0] I_filtered_10b[58] = 013;
    reg [9:0] I_filtered_10b[57] = 016;
    reg [9:0] I_filtered_10b[56] = 018;
    reg [9:0] I_filtered_10b[55] = 01C;
    reg [9:0] I_filtered_10b[54] = 020;
    reg [9:0] I_filtered_10b[53] = 024;
    reg [9:0] I_filtered_10b[52] = 029;
    reg [9:0] I_filtered_10b[51] = 02D;
    reg [9:0] I_filtered_10b[50] = 030;
    reg [9:0] I_filtered_10b[49] = 02F;
    reg [9:0] I_filtered_10b[48] = 02C;
    reg [9:0] I_filtered_10b[47] = 026;
    reg [9:0] I_filtered_10b[46] = 01B;
    reg [9:0] I_filtered_10b[45] = 00E;
    reg [9:0] I_filtered_10b[44] = 3FD;
    reg [9:0] I_filtered_10b[43] = 3EA;
    reg [9:0] I_filtered_10b[42] = 3D2;
    reg [9:0] I_filtered_10b[41] = 3BC;
    reg [9:0] I_filtered_10b[40] = 3A3;
    reg [9:0] I_filtered_10b[39] = 38D;
    reg [9:0] I_filtered_10b[38] = 37A;
    reg [9:0] I_filtered_10b[37] = 36C;
    reg [9:0] I_filtered_10b[36] = 362;
    reg [9:0] I_filtered_10b[35] = 35E;
    reg [9:0] I_filtered_10b[34] = 360;
    reg [9:0] I_filtered_10b[33] = 368;
    reg [9:0] I_filtered_10b[32] = 375;
    reg [9:0] I_filtered_10b[31] = 385;
    reg [9:0] I_filtered_10b[30] = 399;
    reg [9:0] I_filtered_10b[29] = 3AF;
    reg [9:0] I_filtered_10b[28] = 3C4;
    reg [9:0] I_filtered_10b[27] = 3D9;
    reg [9:0] I_filtered_10b[26] = 3EA;
    reg [9:0] I_filtered_10b[25] = 3F8;
    reg [9:0] I_filtered_10b[24] = 003;
    reg [9:0] I_filtered_10b[23] = 00C;
    reg [9:0] I_filtered_10b[22] = 00F;
    reg [9:0] I_filtered_10b[21] = 010;
    reg [9:0] I_filtered_10b[20] = 010;
    reg [9:0] I_filtered_10b[19] = 00D;
    reg [9:0] I_filtered_10b[18] = 009;
    reg [9:0] I_filtered_10b[17] = 006;
    reg [9:0] I_filtered_10b[16] = 002;
    reg [9:0] I_filtered_10b[15] = 3FF;
    reg [9:0] I_filtered_10b[14] = 3FE;
    reg [9:0] I_filtered_10b[13] = 3FC;
    reg [9:0] I_filtered_10b[12] = 3FC;
    reg [9:0] I_filtered_10b[11] = 3FC;
    reg [9:0] I_filtered_10b[10] = 3FE;
    reg [9:0] I_filtered_10b[9] = 000;
    reg [9:0] I_filtered_10b[8] = 001;
    reg [9:0] I_filtered_10b[7] = 002;
    reg [9:0] I_filtered_10b[6] = 002;
    reg [9:0] I_filtered_10b[5] = 004;
    reg [9:0] I_filtered_10b[4] = 002;
    reg [9:0] I_filtered_10b[3] = 002;
    reg [9:0] I_filtered_10b[2] = 001;
    reg [9:0] I_filtered_10b[1] = 000;
    reg [9:0] I_filtered_10b[0] = 000;


    // Q Channel 10b Expected output
    reg [9:0] Q_filtered_10b[1733] = 000;
    reg [9:0] Q_filtered_10b[1732] = 000;
    reg [9:0] Q_filtered_10b[1731] = 000;
    reg [9:0] Q_filtered_10b[1730] = 000;
    reg [9:0] Q_filtered_10b[1729] = 000;
    reg [9:0] Q_filtered_10b[1728] = 000;
    reg [9:0] Q_filtered_10b[1727] = 000;
    reg [9:0] Q_filtered_10b[1726] = 000;
    reg [9:0] Q_filtered_10b[1725] = 000;
    reg [9:0] Q_filtered_10b[1724] = 000;
    reg [9:0] Q_filtered_10b[1723] = 000;
    reg [9:0] Q_filtered_10b[1722] = 000;
    reg [9:0] Q_filtered_10b[1721] = 000;
    reg [9:0] Q_filtered_10b[1720] = 000;
    reg [9:0] Q_filtered_10b[1719] = 001;
    reg [9:0] Q_filtered_10b[1718] = 002;
    reg [9:0] Q_filtered_10b[1717] = 002;
    reg [9:0] Q_filtered_10b[1716] = 004;
    reg [9:0] Q_filtered_10b[1715] = 002;
    reg [9:0] Q_filtered_10b[1714] = 002;
    reg [9:0] Q_filtered_10b[1713] = 001;
    reg [9:0] Q_filtered_10b[1712] = 000;
    reg [9:0] Q_filtered_10b[1711] = 3FE;
    reg [9:0] Q_filtered_10b[1710] = 3FC;
    reg [9:0] Q_filtered_10b[1709] = 3FC;
    reg [9:0] Q_filtered_10b[1708] = 3FC;
    reg [9:0] Q_filtered_10b[1707] = 3FE;
    reg [9:0] Q_filtered_10b[1706] = 3FE;
    reg [9:0] Q_filtered_10b[1705] = 001;
    reg [9:0] Q_filtered_10b[1704] = 005;
    reg [9:0] Q_filtered_10b[1703] = 006;
    reg [9:0] Q_filtered_10b[1702] = 00B;
    reg [9:0] Q_filtered_10b[1701] = 00D;
    reg [9:0] Q_filtered_10b[1700] = 00E;
    reg [9:0] Q_filtered_10b[1699] = 00E;
    reg [9:0] Q_filtered_10b[1698] = 00B;
    reg [9:0] Q_filtered_10b[1697] = 005;
    reg [9:0] Q_filtered_10b[1696] = 3FB;
    reg [9:0] Q_filtered_10b[1695] = 3EE;
    reg [9:0] Q_filtered_10b[1694] = 3DD;
    reg [9:0] Q_filtered_10b[1693] = 3CA;
    reg [9:0] Q_filtered_10b[1692] = 3B4;
    reg [9:0] Q_filtered_10b[1691] = 39F;
    reg [9:0] Q_filtered_10b[1690] = 38C;
    reg [9:0] Q_filtered_10b[1689] = 37C;
    reg [9:0] Q_filtered_10b[1688] = 36F;
    reg [9:0] Q_filtered_10b[1687] = 369;
    reg [9:0] Q_filtered_10b[1686] = 369;
    reg [9:0] Q_filtered_10b[1685] = 36F;
    reg [9:0] Q_filtered_10b[1684] = 37D;
    reg [9:0] Q_filtered_10b[1683] = 38E;
    reg [9:0] Q_filtered_10b[1682] = 3A4;
    reg [9:0] Q_filtered_10b[1681] = 3BD;
    reg [9:0] Q_filtered_10b[1680] = 3D8;
    reg [9:0] Q_filtered_10b[1679] = 3F1;
    reg [9:0] Q_filtered_10b[1678] = 00A;
    reg [9:0] Q_filtered_10b[1677] = 020;
    reg [9:0] Q_filtered_10b[1676] = 033;
    reg [9:0] Q_filtered_10b[1675] = 041;
    reg [9:0] Q_filtered_10b[1674] = 04E;
    reg [9:0] Q_filtered_10b[1673] = 055;
    reg [9:0] Q_filtered_10b[1672] = 05C;
    reg [9:0] Q_filtered_10b[1671] = 060;
    reg [9:0] Q_filtered_10b[1670] = 061;
    reg [9:0] Q_filtered_10b[1669] = 061;
    reg [9:0] Q_filtered_10b[1668] = 064;
    reg [9:0] Q_filtered_10b[1667] = 066;
    reg [9:0] Q_filtered_10b[1666] = 067;
    reg [9:0] Q_filtered_10b[1665] = 06B;
    reg [9:0] Q_filtered_10b[1664] = 06F;
    reg [9:0] Q_filtered_10b[1663] = 071;
    reg [9:0] Q_filtered_10b[1662] = 074;
    reg [9:0] Q_filtered_10b[1661] = 077;
    reg [9:0] Q_filtered_10b[1660] = 078;
    reg [9:0] Q_filtered_10b[1659] = 079;
    reg [9:0] Q_filtered_10b[1658] = 079;
    reg [9:0] Q_filtered_10b[1657] = 079;
    reg [9:0] Q_filtered_10b[1656] = 07A;
    reg [9:0] Q_filtered_10b[1655] = 07C;
    reg [9:0] Q_filtered_10b[1654] = 07D;
    reg [9:0] Q_filtered_10b[1653] = 081;
    reg [9:0] Q_filtered_10b[1652] = 086;
    reg [9:0] Q_filtered_10b[1651] = 088;
    reg [9:0] Q_filtered_10b[1650] = 08F;
    reg [9:0] Q_filtered_10b[1649] = 093;
    reg [9:0] Q_filtered_10b[1648] = 093;
    reg [9:0] Q_filtered_10b[1647] = 08E;
    reg [9:0] Q_filtered_10b[1646] = 089;
    reg [9:0] Q_filtered_10b[1645] = 07A;
    reg [9:0] Q_filtered_10b[1644] = 067;
    reg [9:0] Q_filtered_10b[1643] = 04F;
    reg [9:0] Q_filtered_10b[1642] = 031;
    reg [9:0] Q_filtered_10b[1641] = 011;
    reg [9:0] Q_filtered_10b[1640] = 3F0;
    reg [9:0] Q_filtered_10b[1639] = 3CB;
    reg [9:0] Q_filtered_10b[1638] = 3AC;
    reg [9:0] Q_filtered_10b[1637] = 38D;
    reg [9:0] Q_filtered_10b[1636] = 376;
    reg [9:0] Q_filtered_10b[1635] = 364;
    reg [9:0] Q_filtered_10b[1634] = 35C;
    reg [9:0] Q_filtered_10b[1633] = 359;
    reg [9:0] Q_filtered_10b[1632] = 362;
    reg [9:0] Q_filtered_10b[1631] = 376;
    reg [9:0] Q_filtered_10b[1630] = 38F;
    reg [9:0] Q_filtered_10b[1629] = 3AE;
    reg [9:0] Q_filtered_10b[1628] = 3D1;
    reg [9:0] Q_filtered_10b[1627] = 3F9;
    reg [9:0] Q_filtered_10b[1626] = 01D;
    reg [9:0] Q_filtered_10b[1625] = 03C;
    reg [9:0] Q_filtered_10b[1624] = 057;
    reg [9:0] Q_filtered_10b[1623] = 06B;
    reg [9:0] Q_filtered_10b[1622] = 076;
    reg [9:0] Q_filtered_10b[1621] = 076;
    reg [9:0] Q_filtered_10b[1620] = 071;
    reg [9:0] Q_filtered_10b[1619] = 061;
    reg [9:0] Q_filtered_10b[1618] = 04A;
    reg [9:0] Q_filtered_10b[1617] = 02A;
    reg [9:0] Q_filtered_10b[1616] = 008;
    reg [9:0] Q_filtered_10b[1615] = 3E0;
    reg [9:0] Q_filtered_10b[1614] = 3B7;
    reg [9:0] Q_filtered_10b[1613] = 392;
    reg [9:0] Q_filtered_10b[1612] = 36F;
    reg [9:0] Q_filtered_10b[1611] = 352;
    reg [9:0] Q_filtered_10b[1610] = 33C;
    reg [9:0] Q_filtered_10b[1609] = 32F;
    reg [9:0] Q_filtered_10b[1608] = 32E;
    reg [9:0] Q_filtered_10b[1607] = 331;
    reg [9:0] Q_filtered_10b[1606] = 33F;
    reg [9:0] Q_filtered_10b[1605] = 352;
    reg [9:0] Q_filtered_10b[1604] = 36D;
    reg [9:0] Q_filtered_10b[1603] = 387;
    reg [9:0] Q_filtered_10b[1602] = 3A8;
    reg [9:0] Q_filtered_10b[1601] = 3C8;
    reg [9:0] Q_filtered_10b[1600] = 3E3;
    reg [9:0] Q_filtered_10b[1599] = 3FF;
    reg [9:0] Q_filtered_10b[1598] = 011;
    reg [9:0] Q_filtered_10b[1597] = 021;
    reg [9:0] Q_filtered_10b[1596] = 02A;
    reg [9:0] Q_filtered_10b[1595] = 02D;
    reg [9:0] Q_filtered_10b[1594] = 02B;
    reg [9:0] Q_filtered_10b[1593] = 028;
    reg [9:0] Q_filtered_10b[1592] = 025;
    reg [9:0] Q_filtered_10b[1591] = 01E;
    reg [9:0] Q_filtered_10b[1590] = 01D;
    reg [9:0] Q_filtered_10b[1589] = 01A;
    reg [9:0] Q_filtered_10b[1588] = 01B;
    reg [9:0] Q_filtered_10b[1587] = 01F;
    reg [9:0] Q_filtered_10b[1586] = 021;
    reg [9:0] Q_filtered_10b[1585] = 027;
    reg [9:0] Q_filtered_10b[1584] = 02A;
    reg [9:0] Q_filtered_10b[1583] = 02C;
    reg [9:0] Q_filtered_10b[1582] = 02D;
    reg [9:0] Q_filtered_10b[1581] = 028;
    reg [9:0] Q_filtered_10b[1580] = 01E;
    reg [9:0] Q_filtered_10b[1579] = 00E;
    reg [9:0] Q_filtered_10b[1578] = 3FC;
    reg [9:0] Q_filtered_10b[1577] = 3E1;
    reg [9:0] Q_filtered_10b[1576] = 3C6;
    reg [9:0] Q_filtered_10b[1575] = 3A7;
    reg [9:0] Q_filtered_10b[1574] = 389;
    reg [9:0] Q_filtered_10b[1573] = 36F;
    reg [9:0] Q_filtered_10b[1572] = 359;
    reg [9:0] Q_filtered_10b[1571] = 348;
    reg [9:0] Q_filtered_10b[1570] = 33C;
    reg [9:0] Q_filtered_10b[1569] = 339;
    reg [9:0] Q_filtered_10b[1568] = 33A;
    reg [9:0] Q_filtered_10b[1567] = 343;
    reg [9:0] Q_filtered_10b[1566] = 351;
    reg [9:0] Q_filtered_10b[1565] = 364;
    reg [9:0] Q_filtered_10b[1564] = 378;
    reg [9:0] Q_filtered_10b[1563] = 390;
    reg [9:0] Q_filtered_10b[1562] = 3A7;
    reg [9:0] Q_filtered_10b[1561] = 3BC;
    reg [9:0] Q_filtered_10b[1560] = 3D0;
    reg [9:0] Q_filtered_10b[1559] = 3DD;
    reg [9:0] Q_filtered_10b[1558] = 3E8;
    reg [9:0] Q_filtered_10b[1557] = 3F0;
    reg [9:0] Q_filtered_10b[1556] = 3F4;
    reg [9:0] Q_filtered_10b[1555] = 3F5;
    reg [9:0] Q_filtered_10b[1554] = 3F7;
    reg [9:0] Q_filtered_10b[1553] = 3F8;
    reg [9:0] Q_filtered_10b[1552] = 3F8;
    reg [9:0] Q_filtered_10b[1551] = 3FC;
    reg [9:0] Q_filtered_10b[1550] = 3FD;
    reg [9:0] Q_filtered_10b[1549] = 001;
    reg [9:0] Q_filtered_10b[1548] = 009;
    reg [9:0] Q_filtered_10b[1547] = 00E;
    reg [9:0] Q_filtered_10b[1546] = 017;
    reg [9:0] Q_filtered_10b[1545] = 01C;
    reg [9:0] Q_filtered_10b[1544] = 022;
    reg [9:0] Q_filtered_10b[1543] = 027;
    reg [9:0] Q_filtered_10b[1542] = 029;
    reg [9:0] Q_filtered_10b[1541] = 026;
    reg [9:0] Q_filtered_10b[1540] = 01E;
    reg [9:0] Q_filtered_10b[1539] = 014;
    reg [9:0] Q_filtered_10b[1538] = 004;
    reg [9:0] Q_filtered_10b[1537] = 3F4;
    reg [9:0] Q_filtered_10b[1536] = 3DF;
    reg [9:0] Q_filtered_10b[1535] = 3CA;
    reg [9:0] Q_filtered_10b[1534] = 3BB;
    reg [9:0] Q_filtered_10b[1533] = 3AB;
    reg [9:0] Q_filtered_10b[1532] = 3A0;
    reg [9:0] Q_filtered_10b[1531] = 39A;
    reg [9:0] Q_filtered_10b[1530] = 39A;
    reg [9:0] Q_filtered_10b[1529] = 39E;
    reg [9:0] Q_filtered_10b[1528] = 3AA;
    reg [9:0] Q_filtered_10b[1527] = 3BB;
    reg [9:0] Q_filtered_10b[1526] = 3D2;
    reg [9:0] Q_filtered_10b[1525] = 3EC;
    reg [9:0] Q_filtered_10b[1524] = 009;
    reg [9:0] Q_filtered_10b[1523] = 027;
    reg [9:0] Q_filtered_10b[1522] = 045;
    reg [9:0] Q_filtered_10b[1521] = 05E;
    reg [9:0] Q_filtered_10b[1520] = 077;
    reg [9:0] Q_filtered_10b[1519] = 088;
    reg [9:0] Q_filtered_10b[1518] = 095;
    reg [9:0] Q_filtered_10b[1517] = 099;
    reg [9:0] Q_filtered_10b[1516] = 09A;
    reg [9:0] Q_filtered_10b[1515] = 092;
    reg [9:0] Q_filtered_10b[1514] = 084;
    reg [9:0] Q_filtered_10b[1513] = 070;
    reg [9:0] Q_filtered_10b[1512] = 05A;
    reg [9:0] Q_filtered_10b[1511] = 03F;
    reg [9:0] Q_filtered_10b[1510] = 021;
    reg [9:0] Q_filtered_10b[1509] = 008;
    reg [9:0] Q_filtered_10b[1508] = 3F0;
    reg [9:0] Q_filtered_10b[1507] = 3DE;
    reg [9:0] Q_filtered_10b[1506] = 3CF;
    reg [9:0] Q_filtered_10b[1505] = 3C8;
    reg [9:0] Q_filtered_10b[1504] = 3C8;
    reg [9:0] Q_filtered_10b[1503] = 3CE;
    reg [9:0] Q_filtered_10b[1502] = 3D9;
    reg [9:0] Q_filtered_10b[1501] = 3E8;
    reg [9:0] Q_filtered_10b[1500] = 3FC;
    reg [9:0] Q_filtered_10b[1499] = 010;
    reg [9:0] Q_filtered_10b[1498] = 027;
    reg [9:0] Q_filtered_10b[1497] = 03D;
    reg [9:0] Q_filtered_10b[1496] = 050;
    reg [9:0] Q_filtered_10b[1495] = 062;
    reg [9:0] Q_filtered_10b[1494] = 070;
    reg [9:0] Q_filtered_10b[1493] = 07A;
    reg [9:0] Q_filtered_10b[1492] = 082;
    reg [9:0] Q_filtered_10b[1491] = 083;
    reg [9:0] Q_filtered_10b[1490] = 085;
    reg [9:0] Q_filtered_10b[1489] = 084;
    reg [9:0] Q_filtered_10b[1488] = 083;
    reg [9:0] Q_filtered_10b[1487] = 07E;
    reg [9:0] Q_filtered_10b[1486] = 07F;
    reg [9:0] Q_filtered_10b[1485] = 07D;
    reg [9:0] Q_filtered_10b[1484] = 07D;
    reg [9:0] Q_filtered_10b[1483] = 07E;
    reg [9:0] Q_filtered_10b[1482] = 07E;
    reg [9:0] Q_filtered_10b[1481] = 07F;
    reg [9:0] Q_filtered_10b[1480] = 080;
    reg [9:0] Q_filtered_10b[1479] = 080;
    reg [9:0] Q_filtered_10b[1478] = 07E;
    reg [9:0] Q_filtered_10b[1477] = 07C;
    reg [9:0] Q_filtered_10b[1476] = 076;
    reg [9:0] Q_filtered_10b[1475] = 06F;
    reg [9:0] Q_filtered_10b[1474] = 067;
    reg [9:0] Q_filtered_10b[1473] = 05C;
    reg [9:0] Q_filtered_10b[1472] = 051;
    reg [9:0] Q_filtered_10b[1471] = 046;
    reg [9:0] Q_filtered_10b[1470] = 03A;
    reg [9:0] Q_filtered_10b[1469] = 02E;
    reg [9:0] Q_filtered_10b[1468] = 026;
    reg [9:0] Q_filtered_10b[1467] = 01E;
    reg [9:0] Q_filtered_10b[1466] = 017;
    reg [9:0] Q_filtered_10b[1465] = 011;
    reg [9:0] Q_filtered_10b[1464] = 00E;
    reg [9:0] Q_filtered_10b[1463] = 00A;
    reg [9:0] Q_filtered_10b[1462] = 009;
    reg [9:0] Q_filtered_10b[1461] = 006;
    reg [9:0] Q_filtered_10b[1460] = 003;
    reg [9:0] Q_filtered_10b[1459] = 000;
    reg [9:0] Q_filtered_10b[1458] = 3FD;
    reg [9:0] Q_filtered_10b[1457] = 3F8;
    reg [9:0] Q_filtered_10b[1456] = 3F3;
    reg [9:0] Q_filtered_10b[1455] = 3EC;
    reg [9:0] Q_filtered_10b[1454] = 3E7;
    reg [9:0] Q_filtered_10b[1453] = 3E2;
    reg [9:0] Q_filtered_10b[1452] = 3DE;
    reg [9:0] Q_filtered_10b[1451] = 3DC;
    reg [9:0] Q_filtered_10b[1450] = 3DD;
    reg [9:0] Q_filtered_10b[1449] = 3E2;
    reg [9:0] Q_filtered_10b[1448] = 3E7;
    reg [9:0] Q_filtered_10b[1447] = 3F0;
    reg [9:0] Q_filtered_10b[1446] = 3F8;
    reg [9:0] Q_filtered_10b[1445] = 003;
    reg [9:0] Q_filtered_10b[1444] = 00E;
    reg [9:0] Q_filtered_10b[1443] = 015;
    reg [9:0] Q_filtered_10b[1442] = 01E;
    reg [9:0] Q_filtered_10b[1441] = 023;
    reg [9:0] Q_filtered_10b[1440] = 027;
    reg [9:0] Q_filtered_10b[1439] = 027;
    reg [9:0] Q_filtered_10b[1438] = 026;
    reg [9:0] Q_filtered_10b[1437] = 021;
    reg [9:0] Q_filtered_10b[1436] = 018;
    reg [9:0] Q_filtered_10b[1435] = 00D;
    reg [9:0] Q_filtered_10b[1434] = 3FF;
    reg [9:0] Q_filtered_10b[1433] = 3ED;
    reg [9:0] Q_filtered_10b[1432] = 3DA;
    reg [9:0] Q_filtered_10b[1431] = 3C9;
    reg [9:0] Q_filtered_10b[1430] = 3B8;
    reg [9:0] Q_filtered_10b[1429] = 3AC;
    reg [9:0] Q_filtered_10b[1428] = 3A2;
    reg [9:0] Q_filtered_10b[1427] = 39E;
    reg [9:0] Q_filtered_10b[1426] = 3A0;
    reg [9:0] Q_filtered_10b[1425] = 3A6;
    reg [9:0] Q_filtered_10b[1424] = 3B1;
    reg [9:0] Q_filtered_10b[1423] = 3BE;
    reg [9:0] Q_filtered_10b[1422] = 3D0;
    reg [9:0] Q_filtered_10b[1421] = 3E2;
    reg [9:0] Q_filtered_10b[1420] = 3F5;
    reg [9:0] Q_filtered_10b[1419] = 005;
    reg [9:0] Q_filtered_10b[1418] = 015;
    reg [9:0] Q_filtered_10b[1417] = 024;
    reg [9:0] Q_filtered_10b[1416] = 031;
    reg [9:0] Q_filtered_10b[1415] = 03A;
    reg [9:0] Q_filtered_10b[1414] = 044;
    reg [9:0] Q_filtered_10b[1413] = 04A;
    reg [9:0] Q_filtered_10b[1412] = 053;
    reg [9:0] Q_filtered_10b[1411] = 05A;
    reg [9:0] Q_filtered_10b[1410] = 060;
    reg [9:0] Q_filtered_10b[1409] = 066;
    reg [9:0] Q_filtered_10b[1408] = 070;
    reg [9:0] Q_filtered_10b[1407] = 07B;
    reg [9:0] Q_filtered_10b[1406] = 084;
    reg [9:0] Q_filtered_10b[1405] = 08E;
    reg [9:0] Q_filtered_10b[1404] = 098;
    reg [9:0] Q_filtered_10b[1403] = 09F;
    reg [9:0] Q_filtered_10b[1402] = 0A5;
    reg [9:0] Q_filtered_10b[1401] = 0AA;
    reg [9:0] Q_filtered_10b[1400] = 0AC;
    reg [9:0] Q_filtered_10b[1399] = 0AD;
    reg [9:0] Q_filtered_10b[1398] = 0AC;
    reg [9:0] Q_filtered_10b[1397] = 0AC;
    reg [9:0] Q_filtered_10b[1396] = 0AC;
    reg [9:0] Q_filtered_10b[1395] = 0AE;
    reg [9:0] Q_filtered_10b[1394] = 0B0;
    reg [9:0] Q_filtered_10b[1393] = 0B5;
    reg [9:0] Q_filtered_10b[1392] = 0BB;
    reg [9:0] Q_filtered_10b[1391] = 0BE;
    reg [9:0] Q_filtered_10b[1390] = 0C5;
    reg [9:0] Q_filtered_10b[1389] = 0C9;
    reg [9:0] Q_filtered_10b[1388] = 0C8;
    reg [9:0] Q_filtered_10b[1387] = 0C2;
    reg [9:0] Q_filtered_10b[1386] = 0B9;
    reg [9:0] Q_filtered_10b[1385] = 0A6;
    reg [9:0] Q_filtered_10b[1384] = 090;
    reg [9:0] Q_filtered_10b[1383] = 073;
    reg [9:0] Q_filtered_10b[1382] = 051;
    reg [9:0] Q_filtered_10b[1381] = 02C;
    reg [9:0] Q_filtered_10b[1380] = 008;
    reg [9:0] Q_filtered_10b[1379] = 3E0;
    reg [9:0] Q_filtered_10b[1378] = 3BD;
    reg [9:0] Q_filtered_10b[1377] = 39B;
    reg [9:0] Q_filtered_10b[1376] = 383;
    reg [9:0] Q_filtered_10b[1375] = 36D;
    reg [9:0] Q_filtered_10b[1374] = 361;
    reg [9:0] Q_filtered_10b[1373] = 35B;
    reg [9:0] Q_filtered_10b[1372] = 35D;
    reg [9:0] Q_filtered_10b[1371] = 36A;
    reg [9:0] Q_filtered_10b[1370] = 37A;
    reg [9:0] Q_filtered_10b[1369] = 38E;
    reg [9:0] Q_filtered_10b[1368] = 3A5;
    reg [9:0] Q_filtered_10b[1367] = 3C1;
    reg [9:0] Q_filtered_10b[1366] = 3D7;
    reg [9:0] Q_filtered_10b[1365] = 3EA;
    reg [9:0] Q_filtered_10b[1364] = 3F8;
    reg [9:0] Q_filtered_10b[1363] = 003;
    reg [9:0] Q_filtered_10b[1362] = 007;
    reg [9:0] Q_filtered_10b[1361] = 004;
    reg [9:0] Q_filtered_10b[1360] = 3FE;
    reg [9:0] Q_filtered_10b[1359] = 3F2;
    reg [9:0] Q_filtered_10b[1358] = 3E4;
    reg [9:0] Q_filtered_10b[1357] = 3D0;
    reg [9:0] Q_filtered_10b[1356] = 3BC;
    reg [9:0] Q_filtered_10b[1355] = 3A4;
    reg [9:0] Q_filtered_10b[1354] = 38D;
    reg [9:0] Q_filtered_10b[1353] = 379;
    reg [9:0] Q_filtered_10b[1352] = 365;
    reg [9:0] Q_filtered_10b[1351] = 355;
    reg [9:0] Q_filtered_10b[1350] = 349;
    reg [9:0] Q_filtered_10b[1349] = 342;
    reg [9:0] Q_filtered_10b[1348] = 344;
    reg [9:0] Q_filtered_10b[1347] = 346;
    reg [9:0] Q_filtered_10b[1346] = 34E;
    reg [9:0] Q_filtered_10b[1345] = 357;
    reg [9:0] Q_filtered_10b[1344] = 365;
    reg [9:0] Q_filtered_10b[1343] = 370;
    reg [9:0] Q_filtered_10b[1342] = 37D;
    reg [9:0] Q_filtered_10b[1341] = 387;
    reg [9:0] Q_filtered_10b[1340] = 391;
    reg [9:0] Q_filtered_10b[1339] = 39B;
    reg [9:0] Q_filtered_10b[1338] = 3A2;
    reg [9:0] Q_filtered_10b[1337] = 3A8;
    reg [9:0] Q_filtered_10b[1336] = 3AF;
    reg [9:0] Q_filtered_10b[1335] = 3B6;
    reg [9:0] Q_filtered_10b[1334] = 3BC;
    reg [9:0] Q_filtered_10b[1333] = 3C6;
    reg [9:0] Q_filtered_10b[1332] = 3CF;
    reg [9:0] Q_filtered_10b[1331] = 3DB;
    reg [9:0] Q_filtered_10b[1330] = 3EA;
    reg [9:0] Q_filtered_10b[1329] = 3F8;
    reg [9:0] Q_filtered_10b[1328] = 005;
    reg [9:0] Q_filtered_10b[1327] = 016;
    reg [9:0] Q_filtered_10b[1326] = 025;
    reg [9:0] Q_filtered_10b[1325] = 035;
    reg [9:0] Q_filtered_10b[1324] = 040;
    reg [9:0] Q_filtered_10b[1323] = 04C;
    reg [9:0] Q_filtered_10b[1322] = 055;
    reg [9:0] Q_filtered_10b[1321] = 05D;
    reg [9:0] Q_filtered_10b[1320] = 060;
    reg [9:0] Q_filtered_10b[1319] = 05E;
    reg [9:0] Q_filtered_10b[1318] = 05C;
    reg [9:0] Q_filtered_10b[1317] = 057;
    reg [9:0] Q_filtered_10b[1316] = 053;
    reg [9:0] Q_filtered_10b[1315] = 04A;
    reg [9:0] Q_filtered_10b[1314] = 043;
    reg [9:0] Q_filtered_10b[1313] = 03F;
    reg [9:0] Q_filtered_10b[1312] = 03B;
    reg [9:0] Q_filtered_10b[1311] = 038;
    reg [9:0] Q_filtered_10b[1310] = 038;
    reg [9:0] Q_filtered_10b[1309] = 03A;
    reg [9:0] Q_filtered_10b[1308] = 03E;
    reg [9:0] Q_filtered_10b[1307] = 044;
    reg [9:0] Q_filtered_10b[1306] = 04D;
    reg [9:0] Q_filtered_10b[1305] = 059;
    reg [9:0] Q_filtered_10b[1304] = 067;
    reg [9:0] Q_filtered_10b[1303] = 078;
    reg [9:0] Q_filtered_10b[1302] = 08B;
    reg [9:0] Q_filtered_10b[1301] = 09C;
    reg [9:0] Q_filtered_10b[1300] = 0AC;
    reg [9:0] Q_filtered_10b[1299] = 0B8;
    reg [9:0] Q_filtered_10b[1298] = 0C2;
    reg [9:0] Q_filtered_10b[1297] = 0C6;
    reg [9:0] Q_filtered_10b[1296] = 0C2;
    reg [9:0] Q_filtered_10b[1295] = 0BA;
    reg [9:0] Q_filtered_10b[1294] = 0AC;
    reg [9:0] Q_filtered_10b[1293] = 09C;
    reg [9:0] Q_filtered_10b[1292] = 086;
    reg [9:0] Q_filtered_10b[1291] = 070;
    reg [9:0] Q_filtered_10b[1290] = 055;
    reg [9:0] Q_filtered_10b[1289] = 03E;
    reg [9:0] Q_filtered_10b[1288] = 028;
    reg [9:0] Q_filtered_10b[1287] = 011;
    reg [9:0] Q_filtered_10b[1286] = 003;
    reg [9:0] Q_filtered_10b[1285] = 3F7;
    reg [9:0] Q_filtered_10b[1284] = 3EB;
    reg [9:0] Q_filtered_10b[1283] = 3E4;
    reg [9:0] Q_filtered_10b[1282] = 3DF;
    reg [9:0] Q_filtered_10b[1281] = 3D6;
    reg [9:0] Q_filtered_10b[1280] = 3CE;
    reg [9:0] Q_filtered_10b[1279] = 3C4;
    reg [9:0] Q_filtered_10b[1278] = 3B3;
    reg [9:0] Q_filtered_10b[1277] = 3A4;
    reg [9:0] Q_filtered_10b[1276] = 391;
    reg [9:0] Q_filtered_10b[1275] = 379;
    reg [9:0] Q_filtered_10b[1274] = 366;
    reg [9:0] Q_filtered_10b[1273] = 34E;
    reg [9:0] Q_filtered_10b[1272] = 33E;
    reg [9:0] Q_filtered_10b[1271] = 332;
    reg [9:0] Q_filtered_10b[1270] = 32E;
    reg [9:0] Q_filtered_10b[1269] = 32F;
    reg [9:0] Q_filtered_10b[1268] = 33E;
    reg [9:0] Q_filtered_10b[1267] = 357;
    reg [9:0] Q_filtered_10b[1266] = 376;
    reg [9:0] Q_filtered_10b[1265] = 3A0;
    reg [9:0] Q_filtered_10b[1264] = 3CA;
    reg [9:0] Q_filtered_10b[1263] = 3FA;
    reg [9:0] Q_filtered_10b[1262] = 02B;
    reg [9:0] Q_filtered_10b[1261] = 052;
    reg [9:0] Q_filtered_10b[1260] = 078;
    reg [9:0] Q_filtered_10b[1259] = 094;
    reg [9:0] Q_filtered_10b[1258] = 0A8;
    reg [9:0] Q_filtered_10b[1257] = 0AF;
    reg [9:0] Q_filtered_10b[1256] = 0B0;
    reg [9:0] Q_filtered_10b[1255] = 0A3;
    reg [9:0] Q_filtered_10b[1254] = 08A;
    reg [9:0] Q_filtered_10b[1253] = 06A;
    reg [9:0] Q_filtered_10b[1252] = 044;
    reg [9:0] Q_filtered_10b[1251] = 01A;
    reg [9:0] Q_filtered_10b[1250] = 3EB;
    reg [9:0] Q_filtered_10b[1249] = 3BF;
    reg [9:0] Q_filtered_10b[1248] = 39B;
    reg [9:0] Q_filtered_10b[1247] = 379;
    reg [9:0] Q_filtered_10b[1246] = 360;
    reg [9:0] Q_filtered_10b[1245] = 352;
    reg [9:0] Q_filtered_10b[1244] = 351;
    reg [9:0] Q_filtered_10b[1243] = 355;
    reg [9:0] Q_filtered_10b[1242] = 368;
    reg [9:0] Q_filtered_10b[1241] = 383;
    reg [9:0] Q_filtered_10b[1240] = 3A9;
    reg [9:0] Q_filtered_10b[1239] = 3D2;
    reg [9:0] Q_filtered_10b[1238] = 004;
    reg [9:0] Q_filtered_10b[1237] = 039;
    reg [9:0] Q_filtered_10b[1236] = 068;
    reg [9:0] Q_filtered_10b[1235] = 094;
    reg [9:0] Q_filtered_10b[1234] = 0B8;
    reg [9:0] Q_filtered_10b[1233] = 0D4;
    reg [9:0] Q_filtered_10b[1232] = 0E3;
    reg [9:0] Q_filtered_10b[1231] = 0E3;
    reg [9:0] Q_filtered_10b[1230] = 0DA;
    reg [9:0] Q_filtered_10b[1229] = 0C5;
    reg [9:0] Q_filtered_10b[1228] = 0A9;
    reg [9:0] Q_filtered_10b[1227] = 082;
    reg [9:0] Q_filtered_10b[1226] = 05C;
    reg [9:0] Q_filtered_10b[1225] = 02F;
    reg [9:0] Q_filtered_10b[1224] = 005;
    reg [9:0] Q_filtered_10b[1223] = 3DF;
    reg [9:0] Q_filtered_10b[1222] = 3BB;
    reg [9:0] Q_filtered_10b[1221] = 39F;
    reg [9:0] Q_filtered_10b[1220] = 38A;
    reg [9:0] Q_filtered_10b[1219] = 378;
    reg [9:0] Q_filtered_10b[1218] = 372;
    reg [9:0] Q_filtered_10b[1217] = 36C;
    reg [9:0] Q_filtered_10b[1216] = 369;
    reg [9:0] Q_filtered_10b[1215] = 36A;
    reg [9:0] Q_filtered_10b[1214] = 36E;
    reg [9:0] Q_filtered_10b[1213] = 36A;
    reg [9:0] Q_filtered_10b[1212] = 36A;
    reg [9:0] Q_filtered_10b[1211] = 368;
    reg [9:0] Q_filtered_10b[1210] = 362;
    reg [9:0] Q_filtered_10b[1209] = 35E;
    reg [9:0] Q_filtered_10b[1208] = 358;
    reg [9:0] Q_filtered_10b[1207] = 354;
    reg [9:0] Q_filtered_10b[1206] = 350;
    reg [9:0] Q_filtered_10b[1205] = 34F;
    reg [9:0] Q_filtered_10b[1204] = 34F;
    reg [9:0] Q_filtered_10b[1203] = 354;
    reg [9:0] Q_filtered_10b[1202] = 35B;
    reg [9:0] Q_filtered_10b[1201] = 363;
    reg [9:0] Q_filtered_10b[1200] = 36F;
    reg [9:0] Q_filtered_10b[1199] = 37A;
    reg [9:0] Q_filtered_10b[1198] = 385;
    reg [9:0] Q_filtered_10b[1197] = 391;
    reg [9:0] Q_filtered_10b[1196] = 39B;
    reg [9:0] Q_filtered_10b[1195] = 3A1;
    reg [9:0] Q_filtered_10b[1194] = 3A7;
    reg [9:0] Q_filtered_10b[1193] = 3AE;
    reg [9:0] Q_filtered_10b[1192] = 3B6;
    reg [9:0] Q_filtered_10b[1191] = 3BB;
    reg [9:0] Q_filtered_10b[1190] = 3C5;
    reg [9:0] Q_filtered_10b[1189] = 3CE;
    reg [9:0] Q_filtered_10b[1188] = 3DB;
    reg [9:0] Q_filtered_10b[1187] = 3EA;
    reg [9:0] Q_filtered_10b[1186] = 3FB;
    reg [9:0] Q_filtered_10b[1185] = 00D;
    reg [9:0] Q_filtered_10b[1184] = 020;
    reg [9:0] Q_filtered_10b[1183] = 033;
    reg [9:0] Q_filtered_10b[1182] = 044;
    reg [9:0] Q_filtered_10b[1181] = 051;
    reg [9:0] Q_filtered_10b[1180] = 05B;
    reg [9:0] Q_filtered_10b[1179] = 060;
    reg [9:0] Q_filtered_10b[1178] = 060;
    reg [9:0] Q_filtered_10b[1177] = 05B;
    reg [9:0] Q_filtered_10b[1176] = 051;
    reg [9:0] Q_filtered_10b[1175] = 045;
    reg [9:0] Q_filtered_10b[1174] = 035;
    reg [9:0] Q_filtered_10b[1173] = 024;
    reg [9:0] Q_filtered_10b[1172] = 012;
    reg [9:0] Q_filtered_10b[1171] = 003;
    reg [9:0] Q_filtered_10b[1170] = 3F6;
    reg [9:0] Q_filtered_10b[1169] = 3EF;
    reg [9:0] Q_filtered_10b[1168] = 3E8;
    reg [9:0] Q_filtered_10b[1167] = 3E4;
    reg [9:0] Q_filtered_10b[1166] = 3E4;
    reg [9:0] Q_filtered_10b[1165] = 3E4;
    reg [9:0] Q_filtered_10b[1164] = 3E3;
    reg [9:0] Q_filtered_10b[1163] = 3E1;
    reg [9:0] Q_filtered_10b[1162] = 3DF;
    reg [9:0] Q_filtered_10b[1161] = 3D8;
    reg [9:0] Q_filtered_10b[1160] = 3D2;
    reg [9:0] Q_filtered_10b[1159] = 3C7;
    reg [9:0] Q_filtered_10b[1158] = 3BC;
    reg [9:0] Q_filtered_10b[1157] = 3B3;
    reg [9:0] Q_filtered_10b[1156] = 3A9;
    reg [9:0] Q_filtered_10b[1155] = 3A2;
    reg [9:0] Q_filtered_10b[1154] = 39F;
    reg [9:0] Q_filtered_10b[1153] = 3A0;
    reg [9:0] Q_filtered_10b[1152] = 3A5;
    reg [9:0] Q_filtered_10b[1151] = 3B1;
    reg [9:0] Q_filtered_10b[1150] = 3C1;
    reg [9:0] Q_filtered_10b[1149] = 3D5;
    reg [9:0] Q_filtered_10b[1148] = 3EF;
    reg [9:0] Q_filtered_10b[1147] = 00B;
    reg [9:0] Q_filtered_10b[1146] = 028;
    reg [9:0] Q_filtered_10b[1145] = 044;
    reg [9:0] Q_filtered_10b[1144] = 05D;
    reg [9:0] Q_filtered_10b[1143] = 070;
    reg [9:0] Q_filtered_10b[1142] = 080;
    reg [9:0] Q_filtered_10b[1141] = 08B;
    reg [9:0] Q_filtered_10b[1140] = 08E;
    reg [9:0] Q_filtered_10b[1139] = 08E;
    reg [9:0] Q_filtered_10b[1138] = 08A;
    reg [9:0] Q_filtered_10b[1137] = 083;
    reg [9:0] Q_filtered_10b[1136] = 07A;
    reg [9:0] Q_filtered_10b[1135] = 073;
    reg [9:0] Q_filtered_10b[1134] = 068;
    reg [9:0] Q_filtered_10b[1133] = 060;
    reg [9:0] Q_filtered_10b[1132] = 05C;
    reg [9:0] Q_filtered_10b[1131] = 056;
    reg [9:0] Q_filtered_10b[1130] = 058;
    reg [9:0] Q_filtered_10b[1129] = 057;
    reg [9:0] Q_filtered_10b[1128] = 056;
    reg [9:0] Q_filtered_10b[1127] = 055;
    reg [9:0] Q_filtered_10b[1126] = 054;
    reg [9:0] Q_filtered_10b[1125] = 04A;
    reg [9:0] Q_filtered_10b[1124] = 03C;
    reg [9:0] Q_filtered_10b[1123] = 02B;
    reg [9:0] Q_filtered_10b[1122] = 011;
    reg [9:0] Q_filtered_10b[1121] = 3F8;
    reg [9:0] Q_filtered_10b[1120] = 3DA;
    reg [9:0] Q_filtered_10b[1119] = 3B8;
    reg [9:0] Q_filtered_10b[1118] = 39D;
    reg [9:0] Q_filtered_10b[1117] = 380;
    reg [9:0] Q_filtered_10b[1116] = 36B;
    reg [9:0] Q_filtered_10b[1115] = 35C;
    reg [9:0] Q_filtered_10b[1114] = 356;
    reg [9:0] Q_filtered_10b[1113] = 357;
    reg [9:0] Q_filtered_10b[1112] = 366;
    reg [9:0] Q_filtered_10b[1111] = 381;
    reg [9:0] Q_filtered_10b[1110] = 3A2;
    reg [9:0] Q_filtered_10b[1109] = 3CE;
    reg [9:0] Q_filtered_10b[1108] = 3FB;
    reg [9:0] Q_filtered_10b[1107] = 02F;
    reg [9:0] Q_filtered_10b[1106] = 062;
    reg [9:0] Q_filtered_10b[1105] = 08C;
    reg [9:0] Q_filtered_10b[1104] = 0B4;
    reg [9:0] Q_filtered_10b[1103] = 0D1;
    reg [9:0] Q_filtered_10b[1102] = 0E4;
    reg [9:0] Q_filtered_10b[1101] = 0E8;
    reg [9:0] Q_filtered_10b[1100] = 0E5;
    reg [9:0] Q_filtered_10b[1099] = 0D1;
    reg [9:0] Q_filtered_10b[1098] = 0B1;
    reg [9:0] Q_filtered_10b[1097] = 086;
    reg [9:0] Q_filtered_10b[1096] = 055;
    reg [9:0] Q_filtered_10b[1095] = 01F;
    reg [9:0] Q_filtered_10b[1094] = 3E4;
    reg [9:0] Q_filtered_10b[1093] = 3AB;
    reg [9:0] Q_filtered_10b[1092] = 37B;
    reg [9:0] Q_filtered_10b[1091] = 34D;
    reg [9:0] Q_filtered_10b[1090] = 32C;
    reg [9:0] Q_filtered_10b[1089] = 317;
    reg [9:0] Q_filtered_10b[1088] = 312;
    reg [9:0] Q_filtered_10b[1087] = 315;
    reg [9:0] Q_filtered_10b[1086] = 32A;
    reg [9:0] Q_filtered_10b[1085] = 34B;
    reg [9:0] Q_filtered_10b[1084] = 378;
    reg [9:0] Q_filtered_10b[1083] = 3A9;
    reg [9:0] Q_filtered_10b[1082] = 3E4;
    reg [9:0] Q_filtered_10b[1081] = 023;
    reg [9:0] Q_filtered_10b[1080] = 05C;
    reg [9:0] Q_filtered_10b[1079] = 090;
    reg [9:0] Q_filtered_10b[1078] = 0BA;
    reg [9:0] Q_filtered_10b[1077] = 0DB;
    reg [9:0] Q_filtered_10b[1076] = 0ED;
    reg [9:0] Q_filtered_10b[1075] = 0EE;
    reg [9:0] Q_filtered_10b[1074] = 0E4;
    reg [9:0] Q_filtered_10b[1073] = 0CC;
    reg [9:0] Q_filtered_10b[1072] = 0AB;
    reg [9:0] Q_filtered_10b[1071] = 07E;
    reg [9:0] Q_filtered_10b[1070] = 050;
    reg [9:0] Q_filtered_10b[1069] = 01B;
    reg [9:0] Q_filtered_10b[1068] = 3E8;
    reg [9:0] Q_filtered_10b[1067] = 3B9;
    reg [9:0] Q_filtered_10b[1066] = 38E;
    reg [9:0] Q_filtered_10b[1065] = 36A;
    reg [9:0] Q_filtered_10b[1064] = 34F;
    reg [9:0] Q_filtered_10b[1063] = 33A;
    reg [9:0] Q_filtered_10b[1062] = 333;
    reg [9:0] Q_filtered_10b[1061] = 32E;
    reg [9:0] Q_filtered_10b[1060] = 331;
    reg [9:0] Q_filtered_10b[1059] = 33A;
    reg [9:0] Q_filtered_10b[1058] = 349;
    reg [9:0] Q_filtered_10b[1057] = 353;
    reg [9:0] Q_filtered_10b[1056] = 363;
    reg [9:0] Q_filtered_10b[1055] = 374;
    reg [9:0] Q_filtered_10b[1054] = 37F;
    reg [9:0] Q_filtered_10b[1053] = 38B;
    reg [9:0] Q_filtered_10b[1052] = 392;
    reg [9:0] Q_filtered_10b[1051] = 399;
    reg [9:0] Q_filtered_10b[1050] = 39A;
    reg [9:0] Q_filtered_10b[1049] = 398;
    reg [9:0] Q_filtered_10b[1048] = 394;
    reg [9:0] Q_filtered_10b[1047] = 38F;
    reg [9:0] Q_filtered_10b[1046] = 388;
    reg [9:0] Q_filtered_10b[1045] = 37F;
    reg [9:0] Q_filtered_10b[1044] = 377;
    reg [9:0] Q_filtered_10b[1043] = 36A;
    reg [9:0] Q_filtered_10b[1042] = 35E;
    reg [9:0] Q_filtered_10b[1041] = 356;
    reg [9:0] Q_filtered_10b[1040] = 34D;
    reg [9:0] Q_filtered_10b[1039] = 347;
    reg [9:0] Q_filtered_10b[1038] = 342;
    reg [9:0] Q_filtered_10b[1037] = 342;
    reg [9:0] Q_filtered_10b[1036] = 349;
    reg [9:0] Q_filtered_10b[1035] = 351;
    reg [9:0] Q_filtered_10b[1034] = 35D;
    reg [9:0] Q_filtered_10b[1033] = 368;
    reg [9:0] Q_filtered_10b[1032] = 379;
    reg [9:0] Q_filtered_10b[1031] = 386;
    reg [9:0] Q_filtered_10b[1030] = 398;
    reg [9:0] Q_filtered_10b[1029] = 3A5;
    reg [9:0] Q_filtered_10b[1028] = 3B1;
    reg [9:0] Q_filtered_10b[1027] = 3C1;
    reg [9:0] Q_filtered_10b[1026] = 3C9;
    reg [9:0] Q_filtered_10b[1025] = 3D2;
    reg [9:0] Q_filtered_10b[1024] = 3DB;
    reg [9:0] Q_filtered_10b[1023] = 3E4;
    reg [9:0] Q_filtered_10b[1022] = 3EB;
    reg [9:0] Q_filtered_10b[1021] = 3F7;
    reg [9:0] Q_filtered_10b[1020] = 004;
    reg [9:0] Q_filtered_10b[1019] = 014;
    reg [9:0] Q_filtered_10b[1018] = 02A;
    reg [9:0] Q_filtered_10b[1017] = 043;
    reg [9:0] Q_filtered_10b[1016] = 05E;
    reg [9:0] Q_filtered_10b[1015] = 07B;
    reg [9:0] Q_filtered_10b[1014] = 096;
    reg [9:0] Q_filtered_10b[1013] = 0AF;
    reg [9:0] Q_filtered_10b[1012] = 0C2;
    reg [9:0] Q_filtered_10b[1011] = 0CE;
    reg [9:0] Q_filtered_10b[1010] = 0D2;
    reg [9:0] Q_filtered_10b[1009] = 0CE;
    reg [9:0] Q_filtered_10b[1008] = 0BF;
    reg [9:0] Q_filtered_10b[1007] = 0A9;
    reg [9:0] Q_filtered_10b[1006] = 08E;
    reg [9:0] Q_filtered_10b[1005] = 06C;
    reg [9:0] Q_filtered_10b[1004] = 049;
    reg [9:0] Q_filtered_10b[1003] = 025;
    reg [9:0] Q_filtered_10b[1002] = 003;
    reg [9:0] Q_filtered_10b[1001] = 3E6;
    reg [9:0] Q_filtered_10b[1000] = 3CE;
    reg [9:0] Q_filtered_10b[999] = 3BC;
    reg [9:0] Q_filtered_10b[998] = 3AD;
    reg [9:0] Q_filtered_10b[997] = 3A5;
    reg [9:0] Q_filtered_10b[996] = 39F;
    reg [9:0] Q_filtered_10b[995] = 39C;
    reg [9:0] Q_filtered_10b[994] = 39C;
    reg [9:0] Q_filtered_10b[993] = 39E;
    reg [9:0] Q_filtered_10b[992] = 39B;
    reg [9:0] Q_filtered_10b[991] = 39A;
    reg [9:0] Q_filtered_10b[990] = 398;
    reg [9:0] Q_filtered_10b[989] = 394;
    reg [9:0] Q_filtered_10b[988] = 38F;
    reg [9:0] Q_filtered_10b[987] = 38B;
    reg [9:0] Q_filtered_10b[986] = 388;
    reg [9:0] Q_filtered_10b[985] = 384;
    reg [9:0] Q_filtered_10b[984] = 382;
    reg [9:0] Q_filtered_10b[983] = 383;
    reg [9:0] Q_filtered_10b[982] = 385;
    reg [9:0] Q_filtered_10b[981] = 389;
    reg [9:0] Q_filtered_10b[980] = 38C;
    reg [9:0] Q_filtered_10b[979] = 392;
    reg [9:0] Q_filtered_10b[978] = 397;
    reg [9:0] Q_filtered_10b[977] = 39B;
    reg [9:0] Q_filtered_10b[976] = 39F;
    reg [9:0] Q_filtered_10b[975] = 3A3;
    reg [9:0] Q_filtered_10b[974] = 3A2;
    reg [9:0] Q_filtered_10b[973] = 3A3;
    reg [9:0] Q_filtered_10b[972] = 3A6;
    reg [9:0] Q_filtered_10b[971] = 3AB;
    reg [9:0] Q_filtered_10b[970] = 3B0;
    reg [9:0] Q_filtered_10b[969] = 3BC;
    reg [9:0] Q_filtered_10b[968] = 3CA;
    reg [9:0] Q_filtered_10b[967] = 3DC;
    reg [9:0] Q_filtered_10b[966] = 3F4;
    reg [9:0] Q_filtered_10b[965] = 00D;
    reg [9:0] Q_filtered_10b[964] = 028;
    reg [9:0] Q_filtered_10b[963] = 045;
    reg [9:0] Q_filtered_10b[962] = 05F;
    reg [9:0] Q_filtered_10b[961] = 078;
    reg [9:0] Q_filtered_10b[960] = 08B;
    reg [9:0] Q_filtered_10b[959] = 099;
    reg [9:0] Q_filtered_10b[958] = 09F;
    reg [9:0] Q_filtered_10b[957] = 09F;
    reg [9:0] Q_filtered_10b[956] = 095;
    reg [9:0] Q_filtered_10b[955] = 082;
    reg [9:0] Q_filtered_10b[954] = 06B;
    reg [9:0] Q_filtered_10b[953] = 04D;
    reg [9:0] Q_filtered_10b[952] = 02B;
    reg [9:0] Q_filtered_10b[951] = 006;
    reg [9:0] Q_filtered_10b[950] = 3E5;
    reg [9:0] Q_filtered_10b[949] = 3C7;
    reg [9:0] Q_filtered_10b[948] = 3B1;
    reg [9:0] Q_filtered_10b[947] = 39F;
    reg [9:0] Q_filtered_10b[946] = 395;
    reg [9:0] Q_filtered_10b[945] = 395;
    reg [9:0] Q_filtered_10b[944] = 39B;
    reg [9:0] Q_filtered_10b[943] = 3A6;
    reg [9:0] Q_filtered_10b[942] = 3B5;
    reg [9:0] Q_filtered_10b[941] = 3CA;
    reg [9:0] Q_filtered_10b[940] = 3DE;
    reg [9:0] Q_filtered_10b[939] = 3F5;
    reg [9:0] Q_filtered_10b[938] = 009;
    reg [9:0] Q_filtered_10b[937] = 01A;
    reg [9:0] Q_filtered_10b[936] = 02B;
    reg [9:0] Q_filtered_10b[935] = 037;
    reg [9:0] Q_filtered_10b[934] = 040;
    reg [9:0] Q_filtered_10b[933] = 048;
    reg [9:0] Q_filtered_10b[932] = 04A;
    reg [9:0] Q_filtered_10b[931] = 04F;
    reg [9:0] Q_filtered_10b[930] = 054;
    reg [9:0] Q_filtered_10b[929] = 05A;
    reg [9:0] Q_filtered_10b[928] = 05F;
    reg [9:0] Q_filtered_10b[927] = 06B;
    reg [9:0] Q_filtered_10b[926] = 077;
    reg [9:0] Q_filtered_10b[925] = 085;
    reg [9:0] Q_filtered_10b[924] = 094;
    reg [9:0] Q_filtered_10b[923] = 0A1;
    reg [9:0] Q_filtered_10b[922] = 0AD;
    reg [9:0] Q_filtered_10b[921] = 0B6;
    reg [9:0] Q_filtered_10b[920] = 0BC;
    reg [9:0] Q_filtered_10b[919] = 0BC;
    reg [9:0] Q_filtered_10b[918] = 0BA;
    reg [9:0] Q_filtered_10b[917] = 0B1;
    reg [9:0] Q_filtered_10b[916] = 0A5;
    reg [9:0] Q_filtered_10b[915] = 095;
    reg [9:0] Q_filtered_10b[914] = 083;
    reg [9:0] Q_filtered_10b[913] = 071;
    reg [9:0] Q_filtered_10b[912] = 05F;
    reg [9:0] Q_filtered_10b[911] = 04D;
    reg [9:0] Q_filtered_10b[910] = 03D;
    reg [9:0] Q_filtered_10b[909] = 02F;
    reg [9:0] Q_filtered_10b[908] = 025;
    reg [9:0] Q_filtered_10b[907] = 01A;
    reg [9:0] Q_filtered_10b[906] = 011;
    reg [9:0] Q_filtered_10b[905] = 00A;
    reg [9:0] Q_filtered_10b[904] = 002;
    reg [9:0] Q_filtered_10b[903] = 3FD;
    reg [9:0] Q_filtered_10b[902] = 3F7;
    reg [9:0] Q_filtered_10b[901] = 3F0;
    reg [9:0] Q_filtered_10b[900] = 3E6;
    reg [9:0] Q_filtered_10b[899] = 3DF;
    reg [9:0] Q_filtered_10b[898] = 3D7;
    reg [9:0] Q_filtered_10b[897] = 3CC;
    reg [9:0] Q_filtered_10b[896] = 3C6;
    reg [9:0] Q_filtered_10b[895] = 3C0;
    reg [9:0] Q_filtered_10b[894] = 3BA;
    reg [9:0] Q_filtered_10b[893] = 3B6;
    reg [9:0] Q_filtered_10b[892] = 3B4;
    reg [9:0] Q_filtered_10b[891] = 3B1;
    reg [9:0] Q_filtered_10b[890] = 3AE;
    reg [9:0] Q_filtered_10b[889] = 3AA;
    reg [9:0] Q_filtered_10b[888] = 3A4;
    reg [9:0] Q_filtered_10b[887] = 39E;
    reg [9:0] Q_filtered_10b[886] = 395;
    reg [9:0] Q_filtered_10b[885] = 389;
    reg [9:0] Q_filtered_10b[884] = 381;
    reg [9:0] Q_filtered_10b[883] = 373;
    reg [9:0] Q_filtered_10b[882] = 36A;
    reg [9:0] Q_filtered_10b[881] = 366;
    reg [9:0] Q_filtered_10b[880] = 367;
    reg [9:0] Q_filtered_10b[879] = 36B;
    reg [9:0] Q_filtered_10b[878] = 37C;
    reg [9:0] Q_filtered_10b[877] = 393;
    reg [9:0] Q_filtered_10b[876] = 3B1;
    reg [9:0] Q_filtered_10b[875] = 3D8;
    reg [9:0] Q_filtered_10b[874] = 004;
    reg [9:0] Q_filtered_10b[873] = 035;
    reg [9:0] Q_filtered_10b[872] = 064;
    reg [9:0] Q_filtered_10b[871] = 08E;
    reg [9:0] Q_filtered_10b[870] = 0B2;
    reg [9:0] Q_filtered_10b[869] = 0CE;
    reg [9:0] Q_filtered_10b[868] = 0DF;
    reg [9:0] Q_filtered_10b[867] = 0E3;
    reg [9:0] Q_filtered_10b[866] = 0DC;
    reg [9:0] Q_filtered_10b[865] = 0C9;
    reg [9:0] Q_filtered_10b[864] = 0AD;
    reg [9:0] Q_filtered_10b[863] = 088;
    reg [9:0] Q_filtered_10b[862] = 060;
    reg [9:0] Q_filtered_10b[861] = 031;
    reg [9:0] Q_filtered_10b[860] = 004;
    reg [9:0] Q_filtered_10b[859] = 3DC;
    reg [9:0] Q_filtered_10b[858] = 3B7;
    reg [9:0] Q_filtered_10b[857] = 39C;
    reg [9:0] Q_filtered_10b[856] = 387;
    reg [9:0] Q_filtered_10b[855] = 377;
    reg [9:0] Q_filtered_10b[854] = 372;
    reg [9:0] Q_filtered_10b[853] = 36F;
    reg [9:0] Q_filtered_10b[852] = 36E;
    reg [9:0] Q_filtered_10b[851] = 36E;
    reg [9:0] Q_filtered_10b[850] = 372;
    reg [9:0] Q_filtered_10b[849] = 36D;
    reg [9:0] Q_filtered_10b[848] = 36A;
    reg [9:0] Q_filtered_10b[847] = 363;
    reg [9:0] Q_filtered_10b[846] = 358;
    reg [9:0] Q_filtered_10b[845] = 350;
    reg [9:0] Q_filtered_10b[844] = 347;
    reg [9:0] Q_filtered_10b[843] = 340;
    reg [9:0] Q_filtered_10b[842] = 33D;
    reg [9:0] Q_filtered_10b[841] = 33E;
    reg [9:0] Q_filtered_10b[840] = 345;
    reg [9:0] Q_filtered_10b[839] = 354;
    reg [9:0] Q_filtered_10b[838] = 367;
    reg [9:0] Q_filtered_10b[837] = 37E;
    reg [9:0] Q_filtered_10b[836] = 39C;
    reg [9:0] Q_filtered_10b[835] = 3BA;
    reg [9:0] Q_filtered_10b[834] = 3D7;
    reg [9:0] Q_filtered_10b[833] = 3F6;
    reg [9:0] Q_filtered_10b[832] = 011;
    reg [9:0] Q_filtered_10b[831] = 027;
    reg [9:0] Q_filtered_10b[830] = 038;
    reg [9:0] Q_filtered_10b[829] = 04A;
    reg [9:0] Q_filtered_10b[828] = 055;
    reg [9:0] Q_filtered_10b[827] = 05F;
    reg [9:0] Q_filtered_10b[826] = 068;
    reg [9:0] Q_filtered_10b[825] = 06C;
    reg [9:0] Q_filtered_10b[824] = 070;
    reg [9:0] Q_filtered_10b[823] = 077;
    reg [9:0] Q_filtered_10b[822] = 07F;
    reg [9:0] Q_filtered_10b[821] = 085;
    reg [9:0] Q_filtered_10b[820] = 08E;
    reg [9:0] Q_filtered_10b[819] = 098;
    reg [9:0] Q_filtered_10b[818] = 0A1;
    reg [9:0] Q_filtered_10b[817] = 0A8;
    reg [9:0] Q_filtered_10b[816] = 0AE;
    reg [9:0] Q_filtered_10b[815] = 0B1;
    reg [9:0] Q_filtered_10b[814] = 0B2;
    reg [9:0] Q_filtered_10b[813] = 0AF;
    reg [9:0] Q_filtered_10b[812] = 0AB;
    reg [9:0] Q_filtered_10b[811] = 0A7;
    reg [9:0] Q_filtered_10b[810] = 0A1;
    reg [9:0] Q_filtered_10b[809] = 09E;
    reg [9:0] Q_filtered_10b[808] = 09C;
    reg [9:0] Q_filtered_10b[807] = 099;
    reg [9:0] Q_filtered_10b[806] = 098;
    reg [9:0] Q_filtered_10b[805] = 097;
    reg [9:0] Q_filtered_10b[804] = 097;
    reg [9:0] Q_filtered_10b[803] = 091;
    reg [9:0] Q_filtered_10b[802] = 089;
    reg [9:0] Q_filtered_10b[801] = 07E;
    reg [9:0] Q_filtered_10b[800] = 06C;
    reg [9:0] Q_filtered_10b[799] = 05B;
    reg [9:0] Q_filtered_10b[798] = 044;
    reg [9:0] Q_filtered_10b[797] = 029;
    reg [9:0] Q_filtered_10b[796] = 00D;
    reg [9:0] Q_filtered_10b[795] = 3F4;
    reg [9:0] Q_filtered_10b[794] = 3D8;
    reg [9:0] Q_filtered_10b[793] = 3BE;
    reg [9:0] Q_filtered_10b[792] = 3A6;
    reg [9:0] Q_filtered_10b[791] = 395;
    reg [9:0] Q_filtered_10b[790] = 383;
    reg [9:0] Q_filtered_10b[789] = 377;
    reg [9:0] Q_filtered_10b[788] = 36E;
    reg [9:0] Q_filtered_10b[787] = 368;
    reg [9:0] Q_filtered_10b[786] = 367;
    reg [9:0] Q_filtered_10b[785] = 367;
    reg [9:0] Q_filtered_10b[784] = 366;
    reg [9:0] Q_filtered_10b[783] = 366;
    reg [9:0] Q_filtered_10b[782] = 369;
    reg [9:0] Q_filtered_10b[781] = 367;
    reg [9:0] Q_filtered_10b[780] = 366;
    reg [9:0] Q_filtered_10b[779] = 360;
    reg [9:0] Q_filtered_10b[778] = 35D;
    reg [9:0] Q_filtered_10b[777] = 357;
    reg [9:0] Q_filtered_10b[776] = 354;
    reg [9:0] Q_filtered_10b[775] = 350;
    reg [9:0] Q_filtered_10b[774] = 350;
    reg [9:0] Q_filtered_10b[773] = 353;
    reg [9:0] Q_filtered_10b[772] = 357;
    reg [9:0] Q_filtered_10b[771] = 35D;
    reg [9:0] Q_filtered_10b[770] = 364;
    reg [9:0] Q_filtered_10b[769] = 36D;
    reg [9:0] Q_filtered_10b[768] = 376;
    reg [9:0] Q_filtered_10b[767] = 37E;
    reg [9:0] Q_filtered_10b[766] = 384;
    reg [9:0] Q_filtered_10b[765] = 38A;
    reg [9:0] Q_filtered_10b[764] = 38E;
    reg [9:0] Q_filtered_10b[763] = 393;
    reg [9:0] Q_filtered_10b[762] = 393;
    reg [9:0] Q_filtered_10b[761] = 394;
    reg [9:0] Q_filtered_10b[760] = 391;
    reg [9:0] Q_filtered_10b[759] = 390;
    reg [9:0] Q_filtered_10b[758] = 38B;
    reg [9:0] Q_filtered_10b[757] = 386;
    reg [9:0] Q_filtered_10b[756] = 37F;
    reg [9:0] Q_filtered_10b[755] = 37C;
    reg [9:0] Q_filtered_10b[754] = 379;
    reg [9:0] Q_filtered_10b[753] = 379;
    reg [9:0] Q_filtered_10b[752] = 378;
    reg [9:0] Q_filtered_10b[751] = 37B;
    reg [9:0] Q_filtered_10b[750] = 382;
    reg [9:0] Q_filtered_10b[749] = 388;
    reg [9:0] Q_filtered_10b[748] = 391;
    reg [9:0] Q_filtered_10b[747] = 398;
    reg [9:0] Q_filtered_10b[746] = 3A2;
    reg [9:0] Q_filtered_10b[745] = 3AA;
    reg [9:0] Q_filtered_10b[744] = 3B5;
    reg [9:0] Q_filtered_10b[743] = 3BB;
    reg [9:0] Q_filtered_10b[742] = 3C2;
    reg [9:0] Q_filtered_10b[741] = 3CC;
    reg [9:0] Q_filtered_10b[740] = 3D1;
    reg [9:0] Q_filtered_10b[739] = 3D7;
    reg [9:0] Q_filtered_10b[738] = 3DD;
    reg [9:0] Q_filtered_10b[737] = 3E4;
    reg [9:0] Q_filtered_10b[736] = 3E9;
    reg [9:0] Q_filtered_10b[735] = 3F2;
    reg [9:0] Q_filtered_10b[734] = 3FC;
    reg [9:0] Q_filtered_10b[733] = 009;
    reg [9:0] Q_filtered_10b[732] = 019;
    reg [9:0] Q_filtered_10b[731] = 02B;
    reg [9:0] Q_filtered_10b[730] = 03E;
    reg [9:0] Q_filtered_10b[729] = 054;
    reg [9:0] Q_filtered_10b[728] = 067;
    reg [9:0] Q_filtered_10b[727] = 07B;
    reg [9:0] Q_filtered_10b[726] = 08A;
    reg [9:0] Q_filtered_10b[725] = 095;
    reg [9:0] Q_filtered_10b[724] = 099;
    reg [9:0] Q_filtered_10b[723] = 099;
    reg [9:0] Q_filtered_10b[722] = 08F;
    reg [9:0] Q_filtered_10b[721] = 07D;
    reg [9:0] Q_filtered_10b[720] = 067;
    reg [9:0] Q_filtered_10b[719] = 04B;
    reg [9:0] Q_filtered_10b[718] = 02A;
    reg [9:0] Q_filtered_10b[717] = 006;
    reg [9:0] Q_filtered_10b[716] = 3E6;
    reg [9:0] Q_filtered_10b[715] = 3C8;
    reg [9:0] Q_filtered_10b[714] = 3B2;
    reg [9:0] Q_filtered_10b[713] = 3A0;
    reg [9:0] Q_filtered_10b[712] = 396;
    reg [9:0] Q_filtered_10b[711] = 395;
    reg [9:0] Q_filtered_10b[710] = 39A;
    reg [9:0] Q_filtered_10b[709] = 3A5;
    reg [9:0] Q_filtered_10b[708] = 3B4;
    reg [9:0] Q_filtered_10b[707] = 3C9;
    reg [9:0] Q_filtered_10b[706] = 3DD;
    reg [9:0] Q_filtered_10b[705] = 3F5;
    reg [9:0] Q_filtered_10b[704] = 00A;
    reg [9:0] Q_filtered_10b[703] = 01B;
    reg [9:0] Q_filtered_10b[702] = 02D;
    reg [9:0] Q_filtered_10b[701] = 038;
    reg [9:0] Q_filtered_10b[700] = 041;
    reg [9:0] Q_filtered_10b[699] = 048;
    reg [9:0] Q_filtered_10b[698] = 04A;
    reg [9:0] Q_filtered_10b[697] = 04E;
    reg [9:0] Q_filtered_10b[696] = 052;
    reg [9:0] Q_filtered_10b[695] = 058;
    reg [9:0] Q_filtered_10b[694] = 05D;
    reg [9:0] Q_filtered_10b[693] = 06A;
    reg [9:0] Q_filtered_10b[692] = 074;
    reg [9:0] Q_filtered_10b[691] = 082;
    reg [9:0] Q_filtered_10b[690] = 093;
    reg [9:0] Q_filtered_10b[689] = 09E;
    reg [9:0] Q_filtered_10b[688] = 0AE;
    reg [9:0] Q_filtered_10b[687] = 0B8;
    reg [9:0] Q_filtered_10b[686] = 0C0;
    reg [9:0] Q_filtered_10b[685] = 0C2;
    reg [9:0] Q_filtered_10b[684] = 0C2;
    reg [9:0] Q_filtered_10b[683] = 0B8;
    reg [9:0] Q_filtered_10b[682] = 0A8;
    reg [9:0] Q_filtered_10b[681] = 093;
    reg [9:0] Q_filtered_10b[680] = 079;
    reg [9:0] Q_filtered_10b[679] = 05A;
    reg [9:0] Q_filtered_10b[678] = 038;
    reg [9:0] Q_filtered_10b[677] = 018;
    reg [9:0] Q_filtered_10b[676] = 3FB;
    reg [9:0] Q_filtered_10b[675] = 3E4;
    reg [9:0] Q_filtered_10b[674] = 3D2;
    reg [9:0] Q_filtered_10b[673] = 3C7;
    reg [9:0] Q_filtered_10b[672] = 3C3;
    reg [9:0] Q_filtered_10b[671] = 3C8;
    reg [9:0] Q_filtered_10b[670] = 3D2;
    reg [9:0] Q_filtered_10b[669] = 3E1;
    reg [9:0] Q_filtered_10b[668] = 3F5;
    reg [9:0] Q_filtered_10b[667] = 00B;
    reg [9:0] Q_filtered_10b[666] = 023;
    reg [9:0] Q_filtered_10b[665] = 03A;
    reg [9:0] Q_filtered_10b[664] = 04D;
    reg [9:0] Q_filtered_10b[663] = 05E;
    reg [9:0] Q_filtered_10b[662] = 06B;
    reg [9:0] Q_filtered_10b[661] = 075;
    reg [9:0] Q_filtered_10b[660] = 07D;
    reg [9:0] Q_filtered_10b[659] = 07E;
    reg [9:0] Q_filtered_10b[658] = 082;
    reg [9:0] Q_filtered_10b[657] = 084;
    reg [9:0] Q_filtered_10b[656] = 086;
    reg [9:0] Q_filtered_10b[655] = 086;
    reg [9:0] Q_filtered_10b[654] = 08D;
    reg [9:0] Q_filtered_10b[653] = 093;
    reg [9:0] Q_filtered_10b[652] = 09A;
    reg [9:0] Q_filtered_10b[651] = 0A2;
    reg [9:0] Q_filtered_10b[650] = 0A8;
    reg [9:0] Q_filtered_10b[649] = 0AD;
    reg [9:0] Q_filtered_10b[648] = 0B1;
    reg [9:0] Q_filtered_10b[647] = 0B3;
    reg [9:0] Q_filtered_10b[646] = 0B1;
    reg [9:0] Q_filtered_10b[645] = 0AE;
    reg [9:0] Q_filtered_10b[644] = 0A7;
    reg [9:0] Q_filtered_10b[643] = 0A0;
    reg [9:0] Q_filtered_10b[642] = 097;
    reg [9:0] Q_filtered_10b[641] = 08D;
    reg [9:0] Q_filtered_10b[640] = 084;
    reg [9:0] Q_filtered_10b[639] = 07D;
    reg [9:0] Q_filtered_10b[638] = 075;
    reg [9:0] Q_filtered_10b[637] = 06D;
    reg [9:0] Q_filtered_10b[636] = 067;
    reg [9:0] Q_filtered_10b[635] = 062;
    reg [9:0] Q_filtered_10b[634] = 059;
    reg [9:0] Q_filtered_10b[633] = 050;
    reg [9:0] Q_filtered_10b[632] = 046;
    reg [9:0] Q_filtered_10b[631] = 037;
    reg [9:0] Q_filtered_10b[630] = 02A;
    reg [9:0] Q_filtered_10b[629] = 019;
    reg [9:0] Q_filtered_10b[628] = 005;
    reg [9:0] Q_filtered_10b[627] = 3EF;
    reg [9:0] Q_filtered_10b[626] = 3DC;
    reg [9:0] Q_filtered_10b[625] = 3C6;
    reg [9:0] Q_filtered_10b[624] = 3B1;
    reg [9:0] Q_filtered_10b[623] = 39D;
    reg [9:0] Q_filtered_10b[622] = 38F;
    reg [9:0] Q_filtered_10b[621] = 380;
    reg [9:0] Q_filtered_10b[620] = 377;
    reg [9:0] Q_filtered_10b[619] = 371;
    reg [9:0] Q_filtered_10b[618] = 36E;
    reg [9:0] Q_filtered_10b[617] = 371;
    reg [9:0] Q_filtered_10b[616] = 374;
    reg [9:0] Q_filtered_10b[615] = 378;
    reg [9:0] Q_filtered_10b[614] = 37C;
    reg [9:0] Q_filtered_10b[613] = 382;
    reg [9:0] Q_filtered_10b[612] = 385;
    reg [9:0] Q_filtered_10b[611] = 387;
    reg [9:0] Q_filtered_10b[610] = 387;
    reg [9:0] Q_filtered_10b[609] = 388;
    reg [9:0] Q_filtered_10b[608] = 387;
    reg [9:0] Q_filtered_10b[607] = 388;
    reg [9:0] Q_filtered_10b[606] = 388;
    reg [9:0] Q_filtered_10b[605] = 38A;
    reg [9:0] Q_filtered_10b[604] = 38D;
    reg [9:0] Q_filtered_10b[603] = 390;
    reg [9:0] Q_filtered_10b[602] = 394;
    reg [9:0] Q_filtered_10b[601] = 398;
    reg [9:0] Q_filtered_10b[600] = 39B;
    reg [9:0] Q_filtered_10b[599] = 3A0;
    reg [9:0] Q_filtered_10b[598] = 3A4;
    reg [9:0] Q_filtered_10b[597] = 3A7;
    reg [9:0] Q_filtered_10b[596] = 3AA;
    reg [9:0] Q_filtered_10b[595] = 3AF;
    reg [9:0] Q_filtered_10b[594] = 3B6;
    reg [9:0] Q_filtered_10b[593] = 3BB;
    reg [9:0] Q_filtered_10b[592] = 3C3;
    reg [9:0] Q_filtered_10b[591] = 3C9;
    reg [9:0] Q_filtered_10b[590] = 3D2;
    reg [9:0] Q_filtered_10b[589] = 3DB;
    reg [9:0] Q_filtered_10b[588] = 3E7;
    reg [9:0] Q_filtered_10b[587] = 3F0;
    reg [9:0] Q_filtered_10b[586] = 3FA;
    reg [9:0] Q_filtered_10b[585] = 006;
    reg [9:0] Q_filtered_10b[584] = 00C;
    reg [9:0] Q_filtered_10b[583] = 013;
    reg [9:0] Q_filtered_10b[582] = 018;
    reg [9:0] Q_filtered_10b[581] = 01C;
    reg [9:0] Q_filtered_10b[580] = 01D;
    reg [9:0] Q_filtered_10b[579] = 01F;
    reg [9:0] Q_filtered_10b[578] = 022;
    reg [9:0] Q_filtered_10b[577] = 025;
    reg [9:0] Q_filtered_10b[576] = 02B;
    reg [9:0] Q_filtered_10b[575] = 032;
    reg [9:0] Q_filtered_10b[574] = 03D;
    reg [9:0] Q_filtered_10b[573] = 048;
    reg [9:0] Q_filtered_10b[572] = 052;
    reg [9:0] Q_filtered_10b[571] = 05D;
    reg [9:0] Q_filtered_10b[570] = 065;
    reg [9:0] Q_filtered_10b[569] = 067;
    reg [9:0] Q_filtered_10b[568] = 066;
    reg [9:0] Q_filtered_10b[567] = 05E;
    reg [9:0] Q_filtered_10b[566] = 04E;
    reg [9:0] Q_filtered_10b[565] = 03A;
    reg [9:0] Q_filtered_10b[564] = 021;
    reg [9:0] Q_filtered_10b[563] = 002;
    reg [9:0] Q_filtered_10b[562] = 3E1;
    reg [9:0] Q_filtered_10b[561] = 3C0;
    reg [9:0] Q_filtered_10b[560] = 39E;
    reg [9:0] Q_filtered_10b[559] = 381;
    reg [9:0] Q_filtered_10b[558] = 368;
    reg [9:0] Q_filtered_10b[557] = 355;
    reg [9:0] Q_filtered_10b[556] = 345;
    reg [9:0] Q_filtered_10b[555] = 33E;
    reg [9:0] Q_filtered_10b[554] = 33A;
    reg [9:0] Q_filtered_10b[553] = 33C;
    reg [9:0] Q_filtered_10b[552] = 343;
    reg [9:0] Q_filtered_10b[551] = 34D;
    reg [9:0] Q_filtered_10b[550] = 356;
    reg [9:0] Q_filtered_10b[549] = 362;
    reg [9:0] Q_filtered_10b[548] = 36F;
    reg [9:0] Q_filtered_10b[547] = 378;
    reg [9:0] Q_filtered_10b[546] = 381;
    reg [9:0] Q_filtered_10b[545] = 385;
    reg [9:0] Q_filtered_10b[544] = 38A;
    reg [9:0] Q_filtered_10b[543] = 38C;
    reg [9:0] Q_filtered_10b[542] = 38D;
    reg [9:0] Q_filtered_10b[541] = 38D;
    reg [9:0] Q_filtered_10b[540] = 38F;
    reg [9:0] Q_filtered_10b[539] = 390;
    reg [9:0] Q_filtered_10b[538] = 392;
    reg [9:0] Q_filtered_10b[537] = 396;
    reg [9:0] Q_filtered_10b[536] = 39A;
    reg [9:0] Q_filtered_10b[535] = 39F;
    reg [9:0] Q_filtered_10b[534] = 3A5;
    reg [9:0] Q_filtered_10b[533] = 3AC;
    reg [9:0] Q_filtered_10b[532] = 3AF;
    reg [9:0] Q_filtered_10b[531] = 3B3;
    reg [9:0] Q_filtered_10b[530] = 3B6;
    reg [9:0] Q_filtered_10b[529] = 3BB;
    reg [9:0] Q_filtered_10b[528] = 3BC;
    reg [9:0] Q_filtered_10b[527] = 3BF;
    reg [9:0] Q_filtered_10b[526] = 3C1;
    reg [9:0] Q_filtered_10b[525] = 3C6;
    reg [9:0] Q_filtered_10b[524] = 3C9;
    reg [9:0] Q_filtered_10b[523] = 3D0;
    reg [9:0] Q_filtered_10b[522] = 3D8;
    reg [9:0] Q_filtered_10b[521] = 3DF;
    reg [9:0] Q_filtered_10b[520] = 3E9;
    reg [9:0] Q_filtered_10b[519] = 3EF;
    reg [9:0] Q_filtered_10b[518] = 3F6;
    reg [9:0] Q_filtered_10b[517] = 3F8;
    reg [9:0] Q_filtered_10b[516] = 3FA;
    reg [9:0] Q_filtered_10b[515] = 3F5;
    reg [9:0] Q_filtered_10b[514] = 3EE;
    reg [9:0] Q_filtered_10b[513] = 3E5;
    reg [9:0] Q_filtered_10b[512] = 3DA;
    reg [9:0] Q_filtered_10b[511] = 3CC;
    reg [9:0] Q_filtered_10b[510] = 3BC;
    reg [9:0] Q_filtered_10b[509] = 3AD;
    reg [9:0] Q_filtered_10b[508] = 3A1;
    reg [9:0] Q_filtered_10b[507] = 395;
    reg [9:0] Q_filtered_10b[506] = 390;
    reg [9:0] Q_filtered_10b[505] = 38A;
    reg [9:0] Q_filtered_10b[504] = 387;
    reg [9:0] Q_filtered_10b[503] = 388;
    reg [9:0] Q_filtered_10b[502] = 388;
    reg [9:0] Q_filtered_10b[501] = 388;
    reg [9:0] Q_filtered_10b[500] = 384;
    reg [9:0] Q_filtered_10b[499] = 382;
    reg [9:0] Q_filtered_10b[498] = 378;
    reg [9:0] Q_filtered_10b[497] = 36F;
    reg [9:0] Q_filtered_10b[496] = 360;
    reg [9:0] Q_filtered_10b[495] = 351;
    reg [9:0] Q_filtered_10b[494] = 346;
    reg [9:0] Q_filtered_10b[493] = 339;
    reg [9:0] Q_filtered_10b[492] = 330;
    reg [9:0] Q_filtered_10b[491] = 32E;
    reg [9:0] Q_filtered_10b[490] = 333;
    reg [9:0] Q_filtered_10b[489] = 33D;
    reg [9:0] Q_filtered_10b[488] = 353;
    reg [9:0] Q_filtered_10b[487] = 36E;
    reg [9:0] Q_filtered_10b[486] = 391;
    reg [9:0] Q_filtered_10b[485] = 3BB;
    reg [9:0] Q_filtered_10b[484] = 3EA;
    reg [9:0] Q_filtered_10b[483] = 018;
    reg [9:0] Q_filtered_10b[482] = 047;
    reg [9:0] Q_filtered_10b[481] = 072;
    reg [9:0] Q_filtered_10b[480] = 096;
    reg [9:0] Q_filtered_10b[479] = 0B2;
    reg [9:0] Q_filtered_10b[478] = 0C8;
    reg [9:0] Q_filtered_10b[477] = 0D2;
    reg [9:0] Q_filtered_10b[476] = 0D5;
    reg [9:0] Q_filtered_10b[475] = 0D0;
    reg [9:0] Q_filtered_10b[474] = 0C3;
    reg [9:0] Q_filtered_10b[473] = 0B2;
    reg [9:0] Q_filtered_10b[472] = 0A0;
    reg [9:0] Q_filtered_10b[471] = 08C;
    reg [9:0] Q_filtered_10b[470] = 077;
    reg [9:0] Q_filtered_10b[469] = 068;
    reg [9:0] Q_filtered_10b[468] = 05A;
    reg [9:0] Q_filtered_10b[467] = 052;
    reg [9:0] Q_filtered_10b[466] = 04B;
    reg [9:0] Q_filtered_10b[465] = 046;
    reg [9:0] Q_filtered_10b[464] = 045;
    reg [9:0] Q_filtered_10b[463] = 043;
    reg [9:0] Q_filtered_10b[462] = 03E;
    reg [9:0] Q_filtered_10b[461] = 039;
    reg [9:0] Q_filtered_10b[460] = 035;
    reg [9:0] Q_filtered_10b[459] = 02A;
    reg [9:0] Q_filtered_10b[458] = 020;
    reg [9:0] Q_filtered_10b[457] = 014;
    reg [9:0] Q_filtered_10b[456] = 007;
    reg [9:0] Q_filtered_10b[455] = 3FB;
    reg [9:0] Q_filtered_10b[454] = 3F2;
    reg [9:0] Q_filtered_10b[453] = 3EB;
    reg [9:0] Q_filtered_10b[452] = 3E4;
    reg [9:0] Q_filtered_10b[451] = 3DE;
    reg [9:0] Q_filtered_10b[450] = 3DD;
    reg [9:0] Q_filtered_10b[449] = 3DC;
    reg [9:0] Q_filtered_10b[448] = 3DD;
    reg [9:0] Q_filtered_10b[447] = 3DE;
    reg [9:0] Q_filtered_10b[446] = 3E1;
    reg [9:0] Q_filtered_10b[445] = 3E2;
    reg [9:0] Q_filtered_10b[444] = 3E4;
    reg [9:0] Q_filtered_10b[443] = 3E4;
    reg [9:0] Q_filtered_10b[442] = 3E3;
    reg [9:0] Q_filtered_10b[441] = 3E0;
    reg [9:0] Q_filtered_10b[440] = 3DF;
    reg [9:0] Q_filtered_10b[439] = 3DE;
    reg [9:0] Q_filtered_10b[438] = 3DE;
    reg [9:0] Q_filtered_10b[437] = 3E1;
    reg [9:0] Q_filtered_10b[436] = 3E6;
    reg [9:0] Q_filtered_10b[435] = 3EE;
    reg [9:0] Q_filtered_10b[434] = 3F7;
    reg [9:0] Q_filtered_10b[433] = 004;
    reg [9:0] Q_filtered_10b[432] = 010;
    reg [9:0] Q_filtered_10b[431] = 01E;
    reg [9:0] Q_filtered_10b[430] = 02C;
    reg [9:0] Q_filtered_10b[429] = 038;
    reg [9:0] Q_filtered_10b[428] = 043;
    reg [9:0] Q_filtered_10b[427] = 04B;
    reg [9:0] Q_filtered_10b[426] = 052;
    reg [9:0] Q_filtered_10b[425] = 055;
    reg [9:0] Q_filtered_10b[424] = 057;
    reg [9:0] Q_filtered_10b[423] = 055;
    reg [9:0] Q_filtered_10b[422] = 050;
    reg [9:0] Q_filtered_10b[421] = 049;
    reg [9:0] Q_filtered_10b[420] = 041;
    reg [9:0] Q_filtered_10b[419] = 039;
    reg [9:0] Q_filtered_10b[418] = 02F;
    reg [9:0] Q_filtered_10b[417] = 025;
    reg [9:0] Q_filtered_10b[416] = 01E;
    reg [9:0] Q_filtered_10b[415] = 016;
    reg [9:0] Q_filtered_10b[414] = 011;
    reg [9:0] Q_filtered_10b[413] = 00D;
    reg [9:0] Q_filtered_10b[412] = 00C;
    reg [9:0] Q_filtered_10b[411] = 00C;
    reg [9:0] Q_filtered_10b[410] = 00E;
    reg [9:0] Q_filtered_10b[409] = 014;
    reg [9:0] Q_filtered_10b[408] = 01B;
    reg [9:0] Q_filtered_10b[407] = 023;
    reg [9:0] Q_filtered_10b[406] = 02D;
    reg [9:0] Q_filtered_10b[405] = 038;
    reg [9:0] Q_filtered_10b[404] = 043;
    reg [9:0] Q_filtered_10b[403] = 04B;
    reg [9:0] Q_filtered_10b[402] = 054;
    reg [9:0] Q_filtered_10b[401] = 05A;
    reg [9:0] Q_filtered_10b[400] = 05D;
    reg [9:0] Q_filtered_10b[399] = 05B;
    reg [9:0] Q_filtered_10b[398] = 057;
    reg [9:0] Q_filtered_10b[397] = 04E;
    reg [9:0] Q_filtered_10b[396] = 042;
    reg [9:0] Q_filtered_10b[395] = 031;
    reg [9:0] Q_filtered_10b[394] = 01F;
    reg [9:0] Q_filtered_10b[393] = 00A;
    reg [9:0] Q_filtered_10b[392] = 3F5;
    reg [9:0] Q_filtered_10b[391] = 3E0;
    reg [9:0] Q_filtered_10b[390] = 3CD;
    reg [9:0] Q_filtered_10b[389] = 3BB;
    reg [9:0] Q_filtered_10b[388] = 3AE;
    reg [9:0] Q_filtered_10b[387] = 3A4;
    reg [9:0] Q_filtered_10b[386] = 3A0;
    reg [9:0] Q_filtered_10b[385] = 39F;
    reg [9:0] Q_filtered_10b[384] = 3A4;
    reg [9:0] Q_filtered_10b[383] = 3AE;
    reg [9:0] Q_filtered_10b[382] = 3BB;
    reg [9:0] Q_filtered_10b[381] = 3CB;
    reg [9:0] Q_filtered_10b[380] = 3DB;
    reg [9:0] Q_filtered_10b[379] = 3ED;
    reg [9:0] Q_filtered_10b[378] = 3FE;
    reg [9:0] Q_filtered_10b[377] = 00C;
    reg [9:0] Q_filtered_10b[376] = 01A;
    reg [9:0] Q_filtered_10b[375] = 024;
    reg [9:0] Q_filtered_10b[374] = 02B;
    reg [9:0] Q_filtered_10b[373] = 02D;
    reg [9:0] Q_filtered_10b[372] = 02E;
    reg [9:0] Q_filtered_10b[371] = 029;
    reg [9:0] Q_filtered_10b[370] = 01F;
    reg [9:0] Q_filtered_10b[369] = 012;
    reg [9:0] Q_filtered_10b[368] = 002;
    reg [9:0] Q_filtered_10b[367] = 3EF;
    reg [9:0] Q_filtered_10b[366] = 3D8;
    reg [9:0] Q_filtered_10b[365] = 3C4;
    reg [9:0] Q_filtered_10b[364] = 3B1;
    reg [9:0] Q_filtered_10b[363] = 3A2;
    reg [9:0] Q_filtered_10b[362] = 396;
    reg [9:0] Q_filtered_10b[361] = 392;
    reg [9:0] Q_filtered_10b[360] = 395;
    reg [9:0] Q_filtered_10b[359] = 39E;
    reg [9:0] Q_filtered_10b[358] = 3AF;
    reg [9:0] Q_filtered_10b[357] = 3C4;
    reg [9:0] Q_filtered_10b[356] = 3E0;
    reg [9:0] Q_filtered_10b[355] = 3FF;
    reg [9:0] Q_filtered_10b[354] = 023;
    reg [9:0] Q_filtered_10b[353] = 045;
    reg [9:0] Q_filtered_10b[352] = 066;
    reg [9:0] Q_filtered_10b[351] = 085;
    reg [9:0] Q_filtered_10b[350] = 09D;
    reg [9:0] Q_filtered_10b[349] = 0B0;
    reg [9:0] Q_filtered_10b[348] = 0BE;
    reg [9:0] Q_filtered_10b[347] = 0C2;
    reg [9:0] Q_filtered_10b[346] = 0C3;
    reg [9:0] Q_filtered_10b[345] = 0BF;
    reg [9:0] Q_filtered_10b[344] = 0B8;
    reg [9:0] Q_filtered_10b[343] = 0AD;
    reg [9:0] Q_filtered_10b[342] = 0A6;
    reg [9:0] Q_filtered_10b[341] = 09D;
    reg [9:0] Q_filtered_10b[340] = 098;
    reg [9:0] Q_filtered_10b[339] = 094;
    reg [9:0] Q_filtered_10b[338] = 090;
    reg [9:0] Q_filtered_10b[337] = 08E;
    reg [9:0] Q_filtered_10b[336] = 08C;
    reg [9:0] Q_filtered_10b[335] = 088;
    reg [9:0] Q_filtered_10b[334] = 083;
    reg [9:0] Q_filtered_10b[333] = 07B;
    reg [9:0] Q_filtered_10b[332] = 06E;
    reg [9:0] Q_filtered_10b[331] = 061;
    reg [9:0] Q_filtered_10b[330] = 050;
    reg [9:0] Q_filtered_10b[329] = 03B;
    reg [9:0] Q_filtered_10b[328] = 026;
    reg [9:0] Q_filtered_10b[327] = 013;
    reg [9:0] Q_filtered_10b[326] = 3FC;
    reg [9:0] Q_filtered_10b[325] = 3E9;
    reg [9:0] Q_filtered_10b[324] = 3D7;
    reg [9:0] Q_filtered_10b[323] = 3CA;
    reg [9:0] Q_filtered_10b[322] = 3BB;
    reg [9:0] Q_filtered_10b[321] = 3B0;
    reg [9:0] Q_filtered_10b[320] = 3A6;
    reg [9:0] Q_filtered_10b[319] = 39D;
    reg [9:0] Q_filtered_10b[318] = 398;
    reg [9:0] Q_filtered_10b[317] = 392;
    reg [9:0] Q_filtered_10b[316] = 38A;
    reg [9:0] Q_filtered_10b[315] = 383;
    reg [9:0] Q_filtered_10b[314] = 37F;
    reg [9:0] Q_filtered_10b[313] = 376;
    reg [9:0] Q_filtered_10b[312] = 36E;
    reg [9:0] Q_filtered_10b[311] = 363;
    reg [9:0] Q_filtered_10b[310] = 35C;
    reg [9:0] Q_filtered_10b[309] = 353;
    reg [9:0] Q_filtered_10b[308] = 34F;
    reg [9:0] Q_filtered_10b[307] = 34A;
    reg [9:0] Q_filtered_10b[306] = 34A;
    reg [9:0] Q_filtered_10b[305] = 34E;
    reg [9:0] Q_filtered_10b[304] = 353;
    reg [9:0] Q_filtered_10b[303] = 35B;
    reg [9:0] Q_filtered_10b[302] = 362;
    reg [9:0] Q_filtered_10b[301] = 36C;
    reg [9:0] Q_filtered_10b[300] = 376;
    reg [9:0] Q_filtered_10b[299] = 37E;
    reg [9:0] Q_filtered_10b[298] = 385;
    reg [9:0] Q_filtered_10b[297] = 38A;
    reg [9:0] Q_filtered_10b[296] = 38E;
    reg [9:0] Q_filtered_10b[295] = 393;
    reg [9:0] Q_filtered_10b[294] = 393;
    reg [9:0] Q_filtered_10b[293] = 394;
    reg [9:0] Q_filtered_10b[292] = 392;
    reg [9:0] Q_filtered_10b[291] = 390;
    reg [9:0] Q_filtered_10b[290] = 38B;
    reg [9:0] Q_filtered_10b[289] = 385;
    reg [9:0] Q_filtered_10b[288] = 37D;
    reg [9:0] Q_filtered_10b[287] = 378;
    reg [9:0] Q_filtered_10b[286] = 374;
    reg [9:0] Q_filtered_10b[285] = 373;
    reg [9:0] Q_filtered_10b[284] = 371;
    reg [9:0] Q_filtered_10b[283] = 375;
    reg [9:0] Q_filtered_10b[282] = 37D;
    reg [9:0] Q_filtered_10b[281] = 385;
    reg [9:0] Q_filtered_10b[280] = 392;
    reg [9:0] Q_filtered_10b[279] = 39C;
    reg [9:0] Q_filtered_10b[278] = 3AC;
    reg [9:0] Q_filtered_10b[277] = 3B9;
    reg [9:0] Q_filtered_10b[276] = 3CB;
    reg [9:0] Q_filtered_10b[275] = 3D8;
    reg [9:0] Q_filtered_10b[274] = 3E5;
    reg [9:0] Q_filtered_10b[273] = 3F5;
    reg [9:0] Q_filtered_10b[272] = 3FE;
    reg [9:0] Q_filtered_10b[271] = 007;
    reg [9:0] Q_filtered_10b[270] = 010;
    reg [9:0] Q_filtered_10b[269] = 017;
    reg [9:0] Q_filtered_10b[268] = 01C;
    reg [9:0] Q_filtered_10b[267] = 025;
    reg [9:0] Q_filtered_10b[266] = 02E;
    reg [9:0] Q_filtered_10b[265] = 03A;
    reg [9:0] Q_filtered_10b[264] = 04B;
    reg [9:0] Q_filtered_10b[263] = 05E;
    reg [9:0] Q_filtered_10b[262] = 074;
    reg [9:0] Q_filtered_10b[261] = 08C;
    reg [9:0] Q_filtered_10b[260] = 0A2;
    reg [9:0] Q_filtered_10b[259] = 0B7;
    reg [9:0] Q_filtered_10b[258] = 0C7;
    reg [9:0] Q_filtered_10b[257] = 0D1;
    reg [9:0] Q_filtered_10b[256] = 0D2;
    reg [9:0] Q_filtered_10b[255] = 0CC;
    reg [9:0] Q_filtered_10b[254] = 0BB;
    reg [9:0] Q_filtered_10b[253] = 0A2;
    reg [9:0] Q_filtered_10b[252] = 082;
    reg [9:0] Q_filtered_10b[251] = 05B;
    reg [9:0] Q_filtered_10b[250] = 032;
    reg [9:0] Q_filtered_10b[249] = 008;
    reg [9:0] Q_filtered_10b[248] = 3DE;
    reg [9:0] Q_filtered_10b[247] = 3BA;
    reg [9:0] Q_filtered_10b[246] = 39B;
    reg [9:0] Q_filtered_10b[245] = 383;
    reg [9:0] Q_filtered_10b[244] = 370;
    reg [9:0] Q_filtered_10b[243] = 367;
    reg [9:0] Q_filtered_10b[242] = 361;
    reg [9:0] Q_filtered_10b[241] = 363;
    reg [9:0] Q_filtered_10b[240] = 36B;
    reg [9:0] Q_filtered_10b[239] = 378;
    reg [9:0] Q_filtered_10b[238] = 383;
    reg [9:0] Q_filtered_10b[237] = 392;
    reg [9:0] Q_filtered_10b[236] = 3A3;
    reg [9:0] Q_filtered_10b[235] = 3AF;
    reg [9:0] Q_filtered_10b[234] = 3BA;
    reg [9:0] Q_filtered_10b[233] = 3C1;
    reg [9:0] Q_filtered_10b[232] = 3C7;
    reg [9:0] Q_filtered_10b[231] = 3C8;
    reg [9:0] Q_filtered_10b[230] = 3C6;
    reg [9:0] Q_filtered_10b[229] = 3C2;
    reg [9:0] Q_filtered_10b[228] = 3BD;
    reg [9:0] Q_filtered_10b[227] = 3B7;
    reg [9:0] Q_filtered_10b[226] = 3AE;
    reg [9:0] Q_filtered_10b[225] = 3A7;
    reg [9:0] Q_filtered_10b[224] = 39E;
    reg [9:0] Q_filtered_10b[223] = 395;
    reg [9:0] Q_filtered_10b[222] = 38E;
    reg [9:0] Q_filtered_10b[221] = 387;
    reg [9:0] Q_filtered_10b[220] = 380;
    reg [9:0] Q_filtered_10b[219] = 37C;
    reg [9:0] Q_filtered_10b[218] = 37A;
    reg [9:0] Q_filtered_10b[217] = 37D;
    reg [9:0] Q_filtered_10b[216] = 37F;
    reg [9:0] Q_filtered_10b[215] = 386;
    reg [9:0] Q_filtered_10b[214] = 38D;
    reg [9:0] Q_filtered_10b[213] = 399;
    reg [9:0] Q_filtered_10b[212] = 3A3;
    reg [9:0] Q_filtered_10b[211] = 3B1;
    reg [9:0] Q_filtered_10b[210] = 3BD;
    reg [9:0] Q_filtered_10b[209] = 3CA;
    reg [9:0] Q_filtered_10b[208] = 3D7;
    reg [9:0] Q_filtered_10b[207] = 3E1;
    reg [9:0] Q_filtered_10b[206] = 3E9;
    reg [9:0] Q_filtered_10b[205] = 3F0;
    reg [9:0] Q_filtered_10b[204] = 3F4;
    reg [9:0] Q_filtered_10b[203] = 3F5;
    reg [9:0] Q_filtered_10b[202] = 3F6;
    reg [9:0] Q_filtered_10b[201] = 3F3;
    reg [9:0] Q_filtered_10b[200] = 3F1;
    reg [9:0] Q_filtered_10b[199] = 3EE;
    reg [9:0] Q_filtered_10b[198] = 3EB;
    reg [9:0] Q_filtered_10b[197] = 3E8;
    reg [9:0] Q_filtered_10b[196] = 3E7;
    reg [9:0] Q_filtered_10b[195] = 3E7;
    reg [9:0] Q_filtered_10b[194] = 3E6;
    reg [9:0] Q_filtered_10b[193] = 3E7;
    reg [9:0] Q_filtered_10b[192] = 3E7;
    reg [9:0] Q_filtered_10b[191] = 3E9;
    reg [9:0] Q_filtered_10b[190] = 3E9;
    reg [9:0] Q_filtered_10b[189] = 3E9;
    reg [9:0] Q_filtered_10b[188] = 3E9;
    reg [9:0] Q_filtered_10b[187] = 3EA;
    reg [9:0] Q_filtered_10b[186] = 3E9;
    reg [9:0] Q_filtered_10b[185] = 3EA;
    reg [9:0] Q_filtered_10b[184] = 3EB;
    reg [9:0] Q_filtered_10b[183] = 3EB;
    reg [9:0] Q_filtered_10b[182] = 3ED;
    reg [9:0] Q_filtered_10b[181] = 3EE;
    reg [9:0] Q_filtered_10b[180] = 3F0;
    reg [9:0] Q_filtered_10b[179] = 3EF;
    reg [9:0] Q_filtered_10b[178] = 3EF;
    reg [9:0] Q_filtered_10b[177] = 3EC;
    reg [9:0] Q_filtered_10b[176] = 3E8;
    reg [9:0] Q_filtered_10b[175] = 3E4;
    reg [9:0] Q_filtered_10b[174] = 3DF;
    reg [9:0] Q_filtered_10b[173] = 3D8;
    reg [9:0] Q_filtered_10b[172] = 3D3;
    reg [9:0] Q_filtered_10b[171] = 3CE;
    reg [9:0] Q_filtered_10b[170] = 3C8;
    reg [9:0] Q_filtered_10b[169] = 3C4;
    reg [9:0] Q_filtered_10b[168] = 3BE;
    reg [9:0] Q_filtered_10b[167] = 3BB;
    reg [9:0] Q_filtered_10b[166] = 3B7;
    reg [9:0] Q_filtered_10b[165] = 3B6;
    reg [9:0] Q_filtered_10b[164] = 3B2;
    reg [9:0] Q_filtered_10b[163] = 3B1;
    reg [9:0] Q_filtered_10b[162] = 3B1;
    reg [9:0] Q_filtered_10b[161] = 3B2;
    reg [9:0] Q_filtered_10b[160] = 3B3;
    reg [9:0] Q_filtered_10b[159] = 3B5;
    reg [9:0] Q_filtered_10b[158] = 3B9;
    reg [9:0] Q_filtered_10b[157] = 3BC;
    reg [9:0] Q_filtered_10b[156] = 3BF;
    reg [9:0] Q_filtered_10b[155] = 3C0;
    reg [9:0] Q_filtered_10b[154] = 3C2;
    reg [9:0] Q_filtered_10b[153] = 3C1;
    reg [9:0] Q_filtered_10b[152] = 3C1;
    reg [9:0] Q_filtered_10b[151] = 3BC;
    reg [9:0] Q_filtered_10b[150] = 3B8;
    reg [9:0] Q_filtered_10b[149] = 3B3;
    reg [9:0] Q_filtered_10b[148] = 3AE;
    reg [9:0] Q_filtered_10b[147] = 3A7;
    reg [9:0] Q_filtered_10b[146] = 39F;
    reg [9:0] Q_filtered_10b[145] = 398;
    reg [9:0] Q_filtered_10b[144] = 392;
    reg [9:0] Q_filtered_10b[143] = 38D;
    reg [9:0] Q_filtered_10b[142] = 38A;
    reg [9:0] Q_filtered_10b[141] = 387;
    reg [9:0] Q_filtered_10b[140] = 386;
    reg [9:0] Q_filtered_10b[139] = 388;
    reg [9:0] Q_filtered_10b[138] = 388;
    reg [9:0] Q_filtered_10b[137] = 38A;
    reg [9:0] Q_filtered_10b[136] = 389;
    reg [9:0] Q_filtered_10b[135] = 38A;
    reg [9:0] Q_filtered_10b[134] = 387;
    reg [9:0] Q_filtered_10b[133] = 385;
    reg [9:0] Q_filtered_10b[132] = 37F;
    reg [9:0] Q_filtered_10b[131] = 37A;
    reg [9:0] Q_filtered_10b[130] = 377;
    reg [9:0] Q_filtered_10b[129] = 373;
    reg [9:0] Q_filtered_10b[128] = 370;
    reg [9:0] Q_filtered_10b[127] = 372;
    reg [9:0] Q_filtered_10b[126] = 377;
    reg [9:0] Q_filtered_10b[125] = 37E;
    reg [9:0] Q_filtered_10b[124] = 38C;
    reg [9:0] Q_filtered_10b[123] = 39A;
    reg [9:0] Q_filtered_10b[122] = 3AE;
    reg [9:0] Q_filtered_10b[121] = 3C4;
    reg [9:0] Q_filtered_10b[120] = 3DE;
    reg [9:0] Q_filtered_10b[119] = 3F6;
    reg [9:0] Q_filtered_10b[118] = 00F;
    reg [9:0] Q_filtered_10b[117] = 027;
    reg [9:0] Q_filtered_10b[116] = 039;
    reg [9:0] Q_filtered_10b[115] = 048;
    reg [9:0] Q_filtered_10b[114] = 054;
    reg [9:0] Q_filtered_10b[113] = 05B;
    reg [9:0] Q_filtered_10b[112] = 05C;
    reg [9:0] Q_filtered_10b[111] = 05C;
    reg [9:0] Q_filtered_10b[110] = 059;
    reg [9:0] Q_filtered_10b[109] = 055;
    reg [9:0] Q_filtered_10b[108] = 053;
    reg [9:0] Q_filtered_10b[107] = 050;
    reg [9:0] Q_filtered_10b[106] = 04F;
    reg [9:0] Q_filtered_10b[105] = 051;
    reg [9:0] Q_filtered_10b[104] = 052;
    reg [9:0] Q_filtered_10b[103] = 057;
    reg [9:0] Q_filtered_10b[102] = 05A;
    reg [9:0] Q_filtered_10b[101] = 05B;
    reg [9:0] Q_filtered_10b[100] = 05B;
    reg [9:0] Q_filtered_10b[99] = 056;
    reg [9:0] Q_filtered_10b[98] = 04B;
    reg [9:0] Q_filtered_10b[97] = 03C;
    reg [9:0] Q_filtered_10b[96] = 02A;
    reg [9:0] Q_filtered_10b[95] = 011;
    reg [9:0] Q_filtered_10b[94] = 3F5;
    reg [9:0] Q_filtered_10b[93] = 3D8;
    reg [9:0] Q_filtered_10b[92] = 3BB;
    reg [9:0] Q_filtered_10b[91] = 3A1;
    reg [9:0] Q_filtered_10b[90] = 38C;
    reg [9:0] Q_filtered_10b[89] = 37C;
    reg [9:0] Q_filtered_10b[88] = 370;
    reg [9:0] Q_filtered_10b[87] = 36C;
    reg [9:0] Q_filtered_10b[86] = 36E;
    reg [9:0] Q_filtered_10b[85] = 374;
    reg [9:0] Q_filtered_10b[84] = 37F;
    reg [9:0] Q_filtered_10b[83] = 38D;
    reg [9:0] Q_filtered_10b[82] = 39B;
    reg [9:0] Q_filtered_10b[81] = 3AA;
    reg [9:0] Q_filtered_10b[80] = 3B7;
    reg [9:0] Q_filtered_10b[79] = 3C2;
    reg [9:0] Q_filtered_10b[78] = 3CC;
    reg [9:0] Q_filtered_10b[77] = 3D3;
    reg [9:0] Q_filtered_10b[76] = 3D9;
    reg [9:0] Q_filtered_10b[75] = 3DF;
    reg [9:0] Q_filtered_10b[74] = 3E4;
    reg [9:0] Q_filtered_10b[73] = 3EB;
    reg [9:0] Q_filtered_10b[72] = 3F4;
    reg [9:0] Q_filtered_10b[71] = 3FE;
    reg [9:0] Q_filtered_10b[70] = 009;
    reg [9:0] Q_filtered_10b[69] = 019;
    reg [9:0] Q_filtered_10b[68] = 02A;
    reg [9:0] Q_filtered_10b[67] = 03A;
    reg [9:0] Q_filtered_10b[66] = 04C;
    reg [9:0] Q_filtered_10b[65] = 05C;
    reg [9:0] Q_filtered_10b[64] = 069;
    reg [9:0] Q_filtered_10b[63] = 074;
    reg [9:0] Q_filtered_10b[62] = 07E;
    reg [9:0] Q_filtered_10b[61] = 083;
    reg [9:0] Q_filtered_10b[60] = 087;
    reg [9:0] Q_filtered_10b[59] = 088;
    reg [9:0] Q_filtered_10b[58] = 086;
    reg [9:0] Q_filtered_10b[57] = 084;
    reg [9:0] Q_filtered_10b[56] = 083;
    reg [9:0] Q_filtered_10b[55] = 081;
    reg [9:0] Q_filtered_10b[54] = 080;
    reg [9:0] Q_filtered_10b[53] = 080;
    reg [9:0] Q_filtered_10b[52] = 080;
    reg [9:0] Q_filtered_10b[51] = 084;
    reg [9:0] Q_filtered_10b[50] = 085;
    reg [9:0] Q_filtered_10b[49] = 086;
    reg [9:0] Q_filtered_10b[48] = 083;
    reg [9:0] Q_filtered_10b[47] = 080;
    reg [9:0] Q_filtered_10b[46] = 078;
    reg [9:0] Q_filtered_10b[45] = 06D;
    reg [9:0] Q_filtered_10b[44] = 05F;
    reg [9:0] Q_filtered_10b[43] = 04E;
    reg [9:0] Q_filtered_10b[42] = 03C;
    reg [9:0] Q_filtered_10b[41] = 029;
    reg [9:0] Q_filtered_10b[40] = 014;
    reg [9:0] Q_filtered_10b[39] = 002;
    reg [9:0] Q_filtered_10b[38] = 3F3;
    reg [9:0] Q_filtered_10b[37] = 3E7;
    reg [9:0] Q_filtered_10b[36] = 3DC;
    reg [9:0] Q_filtered_10b[35] = 3D6;
    reg [9:0] Q_filtered_10b[34] = 3D4;
    reg [9:0] Q_filtered_10b[33] = 3D4;
    reg [9:0] Q_filtered_10b[32] = 3D9;
    reg [9:0] Q_filtered_10b[31] = 3DE;
    reg [9:0] Q_filtered_10b[30] = 3E5;
    reg [9:0] Q_filtered_10b[29] = 3ED;
    reg [9:0] Q_filtered_10b[28] = 3F5;
    reg [9:0] Q_filtered_10b[27] = 3FB;
    reg [9:0] Q_filtered_10b[26] = 000;
    reg [9:0] Q_filtered_10b[25] = 002;
    reg [9:0] Q_filtered_10b[24] = 004;
    reg [9:0] Q_filtered_10b[23] = 004;
    reg [9:0] Q_filtered_10b[22] = 003;
    reg [9:0] Q_filtered_10b[21] = 002;
    reg [9:0] Q_filtered_10b[20] = 000;
    reg [9:0] Q_filtered_10b[19] = 000;
    reg [9:0] Q_filtered_10b[18] = 3FE;
    reg [9:0] Q_filtered_10b[17] = 3FF;
    reg [9:0] Q_filtered_10b[16] = 3FE;
    reg [9:0] Q_filtered_10b[15] = 3FF;
    reg [9:0] Q_filtered_10b[14] = 000;
    reg [9:0] Q_filtered_10b[13] = 3FF;
    reg [9:0] Q_filtered_10b[12] = 3FF;
    reg [9:0] Q_filtered_10b[11] = 3FF;
    reg [9:0] Q_filtered_10b[10] = 000;
    reg [9:0] Q_filtered_10b[9] = 000;
    reg [9:0] Q_filtered_10b[8] = 000;
    reg [9:0] Q_filtered_10b[7] = 000;
    reg [9:0] Q_filtered_10b[6] = 000;
    reg [9:0] Q_filtered_10b[5] = 001;
    reg [9:0] Q_filtered_10b[4] = 000;
    reg [9:0] Q_filtered_10b[3] = 000;
    reg [9:0] Q_filtered_10b[2] = 000;
    reg [9:0] Q_filtered_10b[1] = 000;
    reg [9:0] Q_filtered_10b[0] = 000;


    // I Channel 12b Expected output
    //     first 64 samples only
    reg [11:0] I_filtered_12b[63] = 000;
    reg [11:0] I_filtered_12b[62] = 000;
    reg [11:0] I_filtered_12b[61] = 005;
    reg [11:0] I_filtered_12b[60] = 00A;
    reg [11:0] I_filtered_12b[59] = 00A;
    reg [11:0] I_filtered_12b[58] = 00F;
    reg [11:0] I_filtered_12b[57] = 00A;
    reg [11:0] I_filtered_12b[56] = 00A;
    reg [11:0] I_filtered_12b[55] = 005;
    reg [11:0] I_filtered_12b[54] = 000;
    reg [11:0] I_filtered_12b[53] = FF6;
    reg [11:0] I_filtered_12b[52] = FF1;
    reg [11:0] I_filtered_12b[51] = FF1;
    reg [11:0] I_filtered_12b[50] = FF1;
    reg [11:0] I_filtered_12b[49] = FF6;
    reg [11:0] I_filtered_12b[48] = FFA;
    reg [11:0] I_filtered_12b[47] = 008;
    reg [11:0] I_filtered_12b[46] = 017;
    reg [11:0] I_filtered_12b[45] = 025;
    reg [11:0] I_filtered_12b[44] = 035;
    reg [11:0] I_filtered_12b[43] = 03F;
    reg [11:0] I_filtered_12b[42] = 040;
    reg [11:0] I_filtered_12b[41] = 03C;
    reg [11:0] I_filtered_12b[40] = 02F;
    reg [11:0] I_filtered_12b[39] = 00D;
    reg [11:0] I_filtered_12b[38] = FE0;
    reg [11:0] I_filtered_12b[37] = FA9;
    reg [11:0] I_filtered_12b[36] = F62;
    reg [11:0] I_filtered_12b[35] = F10;
    reg [11:0] I_filtered_12b[34] = EBC;
    reg [11:0] I_filtered_12b[33] = E64;
    reg [11:0] I_filtered_12b[32] = E15;
    reg [11:0] I_filtered_12b[31] = DD2;
    reg [11:0] I_filtered_12b[30] = D9E;
    reg [11:0] I_filtered_12b[29] = D81;
    reg [11:0] I_filtered_12b[28] = D79;
    reg [11:0] I_filtered_12b[27] = D88;
    reg [11:0] I_filtered_12b[26] = DAE;
    reg [11:0] I_filtered_12b[25] = DE9;
    reg [11:0] I_filtered_12b[24] = E35;
    reg [11:0] I_filtered_12b[23] = E8D;
    reg [11:0] I_filtered_12b[22] = EEE;
    reg [11:0] I_filtered_12b[21] = F48;
    reg [11:0] I_filtered_12b[20] = FA6;
    reg [11:0] I_filtered_12b[19] = FF5;
    reg [11:0] I_filtered_12b[18] = 039;
    reg [11:0] I_filtered_12b[17] = 06E;
    reg [11:0] I_filtered_12b[16] = 09A;
    reg [11:0] I_filtered_12b[15] = 0AF;
    reg [11:0] I_filtered_12b[14] = 0BB;
    reg [11:0] I_filtered_12b[13] = 0BF;
    reg [11:0] I_filtered_12b[12] = 0B4;
    reg [11:0] I_filtered_12b[11] = 0A3;
    reg [11:0] I_filtered_12b[10] = 090;
    reg [11:0] I_filtered_12b[9] = 082;
    reg [11:0] I_filtered_12b[8] = 06F;
    reg [11:0] I_filtered_12b[7] = 062;
    reg [11:0] I_filtered_12b[6] = 05A;
    reg [11:0] I_filtered_12b[5] = 04E;
    reg [11:0] I_filtered_12b[4] = 049;
    reg [11:0] I_filtered_12b[3] = 048;
    reg [11:0] I_filtered_12b[2] = 04F;
    reg [11:0] I_filtered_12b[1] = 050;
    reg [11:0] I_filtered_12b[0] = 05F;


    // Q Channel 12b Expected output
    //     first 64 samples only
    reg [11:0] Q_filtered_12b[63] = 000;
    reg [11:0] Q_filtered_12b[62] = 000;
    reg [11:0] Q_filtered_12b[61] = 001;
    reg [11:0] Q_filtered_12b[60] = 002;
    reg [11:0] Q_filtered_12b[59] = 002;
    reg [11:0] Q_filtered_12b[58] = 003;
    reg [11:0] Q_filtered_12b[57] = 002;
    reg [11:0] Q_filtered_12b[56] = 002;
    reg [11:0] Q_filtered_12b[55] = 001;
    reg [11:0] Q_filtered_12b[54] = 000;
    reg [11:0] Q_filtered_12b[53] = FFE;
    reg [11:0] Q_filtered_12b[52] = FFD;
    reg [11:0] Q_filtered_12b[51] = FFD;
    reg [11:0] Q_filtered_12b[50] = FFD;
    reg [11:0] Q_filtered_12b[49] = FFE;
    reg [11:0] Q_filtered_12b[48] = FFA;
    reg [11:0] Q_filtered_12b[47] = FF8;
    reg [11:0] Q_filtered_12b[46] = FFB;
    reg [11:0] Q_filtered_12b[45] = FF8;
    reg [11:0] Q_filtered_12b[44] = 000;
    reg [11:0] Q_filtered_12b[43] = 002;
    reg [11:0] Q_filtered_12b[42] = 007;
    reg [11:0] Q_filtered_12b[41] = 00B;
    reg [11:0] Q_filtered_12b[40] = 012;
    reg [11:0] Q_filtered_12b[39] = 011;
    reg [11:0] Q_filtered_12b[38] = 009;
    reg [11:0] Q_filtered_12b[37] = FFF;
    reg [11:0] Q_filtered_12b[36] = FED;
    reg [11:0] Q_filtered_12b[35] = FD5;
    reg [11:0] Q_filtered_12b[34] = FB2;
    reg [11:0] Q_filtered_12b[33] = F94;
    reg [11:0] Q_filtered_12b[32] = F78;
    reg [11:0] Q_filtered_12b[31] = F62;
    reg [11:0] Q_filtered_12b[30] = F4F;
    reg [11:0] Q_filtered_12b[29] = F4E;
    reg [11:0] Q_filtered_12b[28] = F57;
    reg [11:0] Q_filtered_12b[27] = F71;
    reg [11:0] Q_filtered_12b[26] = F9A;
    reg [11:0] Q_filtered_12b[25] = FCB;
    reg [11:0] Q_filtered_12b[24] = 009;
    reg [11:0] Q_filtered_12b[23] = 052;
    reg [11:0] Q_filtered_12b[22] = 0A3;
    reg [11:0] Q_filtered_12b[21] = 0EF;
    reg [11:0] Q_filtered_12b[20] = 139;
    reg [11:0] Q_filtered_12b[19] = 17E;
    reg [11:0] Q_filtered_12b[18] = 1B4;
    reg [11:0] Q_filtered_12b[17] = 1DF;
    reg [11:0] Q_filtered_12b[16] = 202;
    reg [11:0] Q_filtered_12b[15] = 20E;
    reg [11:0] Q_filtered_12b[14] = 217;
    reg [11:0] Q_filtered_12b[13] = 216;
    reg [11:0] Q_filtered_12b[12] = 20F;
    reg [11:0] Q_filtered_12b[11] = 202;
    reg [11:0] Q_filtered_12b[10] = 201;
    reg [11:0] Q_filtered_12b[9] = 1FF;
    reg [11:0] Q_filtered_12b[8] = 204;
    reg [11:0] Q_filtered_12b[7] = 20B;
    reg [11:0] Q_filtered_12b[6] = 211;
    reg [11:0] Q_filtered_12b[5] = 219;
    reg [11:0] Q_filtered_12b[4] = 220;
    reg [11:0] Q_filtered_12b[3] = 21C;
    reg [11:0] Q_filtered_12b[2] = 20E;
    reg [11:0] Q_filtered_12b[1] = 1F8;
    reg [11:0] Q_filtered_12b[0] = 1D0;
end

endmodule

